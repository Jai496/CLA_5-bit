magic
tech scmos
timestamp 1763383735
<< nwell >>
rect 3209 794 3233 818
rect 3248 808 3282 814
rect 3248 778 3310 808
rect 3276 772 3310 778
rect 3209 739 3233 763
<< ntransistor >>
rect 3220 780 3222 786
rect 3259 731 3261 743
rect 3269 731 3271 743
rect 3287 731 3289 743
rect 3297 731 3299 743
rect 3220 725 3222 731
<< ptransistor >>
rect 3220 800 3222 812
rect 3259 784 3261 808
rect 3269 784 3271 808
rect 3287 778 3289 802
rect 3297 778 3299 802
rect 3220 745 3222 757
<< ndiffusion >>
rect 3219 780 3220 786
rect 3222 780 3223 786
rect 3258 731 3259 743
rect 3261 731 3269 743
rect 3271 731 3272 743
rect 3286 731 3287 743
rect 3289 731 3297 743
rect 3299 731 3300 743
rect 3219 725 3220 731
rect 3222 725 3223 731
<< pdiffusion >>
rect 3219 800 3220 812
rect 3222 800 3223 812
rect 3258 784 3259 808
rect 3261 784 3263 808
rect 3267 784 3269 808
rect 3271 784 3272 808
rect 3286 778 3287 802
rect 3289 778 3291 802
rect 3295 778 3297 802
rect 3299 778 3300 802
rect 3219 745 3220 757
rect 3222 745 3223 757
<< ndcontact >>
rect 3215 780 3219 786
rect 3223 780 3227 786
rect 3254 731 3258 743
rect 3272 731 3276 743
rect 3282 731 3286 743
rect 3300 731 3304 743
rect 3215 725 3219 731
rect 3223 725 3227 731
<< pdcontact >>
rect 3215 800 3219 812
rect 3223 800 3227 812
rect 3254 784 3258 808
rect 3263 784 3267 808
rect 3272 784 3276 808
rect 3282 778 3286 802
rect 3291 778 3295 802
rect 3300 778 3304 802
rect 3215 745 3219 757
rect 3223 745 3227 757
<< polysilicon >>
rect 3220 812 3222 815
rect 3259 808 3261 811
rect 3269 808 3271 811
rect 3220 786 3222 800
rect 3287 802 3289 805
rect 3297 802 3299 805
rect 3220 777 3222 780
rect 3259 775 3261 784
rect 3269 774 3271 784
rect 3220 757 3222 760
rect 3220 731 3222 745
rect 3259 743 3261 770
rect 3269 743 3271 769
rect 3287 767 3289 778
rect 3287 743 3289 763
rect 3297 756 3299 778
rect 3297 743 3299 752
rect 3259 728 3261 731
rect 3269 728 3271 731
rect 3287 728 3289 731
rect 3297 728 3299 731
rect 3220 722 3222 725
<< polycontact >>
rect 3216 789 3220 793
rect 3216 734 3220 738
rect 3285 763 3289 767
rect 3296 752 3300 756
<< metal1 >>
rect 3214 818 3242 821
rect 3215 812 3218 818
rect 3239 817 3242 818
rect 3239 814 3310 817
rect 3182 788 3201 791
rect 3206 789 3216 792
rect 3224 792 3227 800
rect 3254 808 3257 814
rect 3273 808 3276 814
rect 3224 789 3245 792
rect 3224 786 3227 789
rect 3215 776 3218 780
rect 3209 774 3233 776
rect 3209 773 3227 774
rect 3232 773 3233 774
rect 3242 766 3245 789
rect 3283 808 3303 811
rect 3283 802 3286 808
rect 3300 802 3303 808
rect 3264 781 3267 784
rect 3264 778 3282 781
rect 3292 771 3295 778
rect 3292 768 3309 771
rect 3214 765 3233 766
rect 3209 763 3233 765
rect 3242 763 3285 766
rect 3215 757 3218 763
rect 3306 757 3309 768
rect 3271 752 3296 755
rect 3306 753 3313 757
rect 3271 750 3274 752
rect 3182 734 3201 737
rect 3206 734 3216 737
rect 3224 737 3227 745
rect 3236 747 3274 750
rect 3306 749 3309 753
rect 3236 737 3239 747
rect 3277 746 3309 749
rect 3277 743 3280 746
rect 3224 734 3239 737
rect 3224 731 3227 734
rect 3276 740 3282 743
rect 3215 721 3218 725
rect 3236 724 3241 727
rect 3254 727 3257 731
rect 3301 727 3304 731
rect 3246 724 3310 727
rect 3236 721 3239 724
rect 3209 718 3239 721
<< m2contact >>
rect 3201 787 3206 792
rect 3201 733 3206 738
<< pm12contact >>
rect 3257 770 3262 775
rect 3266 769 3271 774
<< metal2 >>
rect 3202 781 3205 787
rect 3202 778 3239 781
rect 3236 775 3239 778
rect 3236 772 3257 775
rect 3266 759 3269 769
rect 3203 756 3269 759
rect 3203 738 3206 756
<< m123contact >>
rect 3209 818 3214 823
rect 3209 765 3214 770
rect 3227 769 3232 774
rect 3241 724 3246 729
<< metal3 >>
rect 3209 770 3212 818
rect 3232 769 3244 772
rect 3241 729 3244 769
<< labels >>
rlabel metal1 3222 764 3225 766 1 vdd
rlabel metal1 3221 818 3224 820 5 vdd
rlabel metal1 3225 774 3226 776 1 gnd
rlabel metal1 3277 724 3280 726 1 gnd
rlabel metal1 3227 718 3231 721 1 gnd
rlabel metal1 3306 753 3313 757 7 out
rlabel metal1 3182 788 3201 791 1 A
rlabel metal1 3182 734 3201 737 1 B
rlabel metal1 3224 789 3245 792 1 A_bar
rlabel metal1 3224 734 3239 737 1 B_bar
<< end >>
