* Static P/G 
* Author: Jai Srikar 2024102041

.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param W_N = 20 * LAMBDA
.param W_P = 2 * W_N

* Inverter (A -> A_bar)
M1 A_bar A VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M2 A_bar A GND GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* Inverter (B -> B_bar)
M3 B_bar B VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M4 B_bar B GND GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* 1. Generate (G) - Static NAND + Inverter (G = A AND B)

* NAND(A, B) -> G_bar
* PUN
M5 G_bar A VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M6 G_bar B VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}

* PDN
M7 G_bar A n_g1 GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}
M8 n_g1 B GND GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* Inverter (G_bar -> G)
M9 G G_bar VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M10 G G_bar GND GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* 2. Propagate (P) - Transmission Gate XOR (P = A XOR B)

* --- XNOR WITH TG ---
* TG1 (passes A when B=1 / B_bar=0)
M11 n_p1 B_bar A VDD CMOSP W={W_P} L={LAMBDA} ; PMOS gate=B_bar
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M12 n_p1 B A GND CMOSN W={W_N} L={LAMBDA}    ; NMOS gate=B
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* TG2 (passes A_bar when B=0 / B_bar=1)
M13 n_p1 B A_bar VDD CMOSP W={W_P} L={LAMBDA} ; PMOS gate=B
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M14 n_p1 B_bar A_bar GND CMOSN W={W_N} L={LAMBDA} ; NMOS gate=B_bar
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}

* --- Output Inverter  ---
M15 P n_p1 VDD VDD CMOSP W={W_P} L={LAMBDA}
+ AS={5*W_P*LAMBDA} PS={10*LAMBDA+2*W_P} AD={5*W_P*LAMBDA} PD={10*LAMBDA+2*W_P}
M16 P n_p1 GND GND CMOSN W={W_N} L={LAMBDA}
+ AS={5*W_N*LAMBDA} PS={10*LAMBDA+2*W_N} AD={5*W_N*LAMBDA} PD={10*LAMBDA+2*W_N}