module dff_tb;
    reg D;
    reg CLK;
    wire Q;

    dff uut (
        .D(D), 
        .CLK(CLK), 
        .Q(Q)
    );

    always #0.5 CLK = ~CLK;

    initial begin
        CLK = 0;
        D = 0;
        $dumpfile("dff_tb.vcd");
        $dumpvars(0, dff_tb);

        #0.25 D = 1;  // Setup for first rising edge (at 1.0ns)
        #1.00 D = 0;  // Hold for first edge, setup for second
        #1.00 D = 1;  // High again
        #2.00 D = 0;
        
        #2.00 $finish;
    end

    initial begin
        $monitor("Time=%t | CLK=%b D=%b | Q=%b", $time, CLK, D, Q);
    end

endmodule