magic
tech scmos
timestamp 1764695306
<< nwell >>
rect -8117 -2648 -8094 -2623
rect -7975 -2651 -7952 -2626
rect -7833 -2649 -7810 -2624
rect -7699 -2642 -7676 -2617
rect -7564 -2648 -7541 -2623
rect -7444 -2647 -7421 -2622
rect -7324 -2647 -7301 -2622
rect -7199 -2646 -7176 -2621
rect -7081 -2646 -7058 -2621
rect -6962 -2644 -6939 -2619
rect -8117 -2691 -8096 -2666
rect -7975 -2694 -7954 -2669
rect -7833 -2692 -7812 -2667
rect -7699 -2685 -7678 -2660
rect -7564 -2691 -7543 -2666
rect -7444 -2690 -7423 -2665
rect -7324 -2690 -7303 -2665
rect -7199 -2689 -7178 -2664
rect -7081 -2689 -7060 -2664
rect -6962 -2687 -6941 -2662
rect -8117 -2733 -8094 -2708
rect -7975 -2736 -7952 -2711
rect -7833 -2734 -7810 -2709
rect -7699 -2727 -7676 -2702
rect -7564 -2733 -7541 -2708
rect -7444 -2732 -7421 -2707
rect -7324 -2732 -7301 -2707
rect -7199 -2731 -7176 -2706
rect -7081 -2731 -7058 -2706
rect -6962 -2729 -6939 -2704
rect -8114 -2821 -8089 -2764
rect -7972 -2824 -7947 -2767
rect -7830 -2822 -7805 -2765
rect -7696 -2815 -7671 -2758
rect -7561 -2821 -7536 -2764
rect -7441 -2820 -7416 -2763
rect -7321 -2820 -7296 -2763
rect -7196 -2819 -7171 -2762
rect -7078 -2819 -7053 -2762
rect -6959 -2817 -6934 -2760
rect -8117 -2864 -8094 -2839
rect -7975 -2867 -7952 -2842
rect -7833 -2865 -7810 -2840
rect -7699 -2858 -7676 -2833
rect -7564 -2864 -7541 -2839
rect -7444 -2863 -7421 -2838
rect -7324 -2863 -7301 -2838
rect -7199 -2862 -7176 -2837
rect -7081 -2862 -7058 -2837
rect -6962 -2860 -6939 -2835
rect -8117 -2907 -8096 -2882
rect -7975 -2910 -7954 -2885
rect -7833 -2908 -7812 -2883
rect -7699 -2901 -7678 -2876
rect -7564 -2907 -7543 -2882
rect -7444 -2906 -7423 -2881
rect -7324 -2906 -7303 -2881
rect -7199 -2905 -7178 -2880
rect -7081 -2905 -7060 -2880
rect -6962 -2903 -6941 -2878
rect -8117 -2949 -8094 -2924
rect -7975 -2952 -7952 -2927
rect -7833 -2950 -7810 -2925
rect -7699 -2943 -7676 -2918
rect -7564 -2949 -7541 -2924
rect -7444 -2948 -7421 -2923
rect -7324 -2948 -7301 -2923
rect -7199 -2947 -7176 -2922
rect -7081 -2947 -7058 -2922
rect -6962 -2945 -6939 -2920
rect -8114 -3037 -8089 -2980
rect -7972 -3040 -7947 -2983
rect -7830 -3038 -7805 -2981
rect -7696 -3031 -7671 -2974
rect -7561 -3037 -7536 -2980
rect -7441 -3036 -7416 -2979
rect -7321 -3036 -7296 -2979
rect -7196 -3035 -7171 -2978
rect -7078 -3035 -7053 -2978
rect -6959 -3033 -6934 -2976
rect -5243 -3036 -5219 -2984
rect -3739 -3211 -3715 -3187
rect -3700 -3197 -3666 -3191
rect -5109 -3273 -5085 -3211
rect -4937 -3274 -4913 -3212
rect -4763 -3274 -4739 -3212
rect -4639 -3275 -4615 -3213
rect -4499 -3278 -4475 -3216
rect -3700 -3227 -3638 -3197
rect -3672 -3233 -3638 -3227
rect -3739 -3266 -3715 -3242
rect -3564 -3248 -3539 -3225
rect -3521 -3248 -3496 -3227
rect -3479 -3248 -3454 -3225
rect -3423 -3245 -3366 -3220
rect -3348 -3248 -3323 -3225
rect -3305 -3248 -3280 -3227
rect -3263 -3248 -3238 -3225
rect -3207 -3245 -3150 -3220
rect -4300 -3395 -4276 -3343
rect -3808 -3395 -3784 -3371
rect -3769 -3381 -3735 -3375
rect -3769 -3411 -3707 -3381
rect -3741 -3417 -3707 -3411
rect -6083 -3470 -6059 -3446
rect -3808 -3450 -3784 -3426
rect -3569 -3432 -3544 -3409
rect -3526 -3432 -3501 -3411
rect -3484 -3432 -3459 -3409
rect -3428 -3429 -3371 -3404
rect -3353 -3432 -3328 -3409
rect -3310 -3432 -3285 -3411
rect -3268 -3432 -3243 -3409
rect -3212 -3429 -3155 -3404
rect -6044 -3456 -6010 -3450
rect -6044 -3486 -5982 -3456
rect -6016 -3492 -5982 -3486
rect -6083 -3525 -6059 -3501
rect -4299 -3526 -4275 -3474
rect -3813 -3525 -3789 -3501
rect -3774 -3511 -3740 -3505
rect -3774 -3541 -3712 -3511
rect -3746 -3547 -3712 -3541
rect -3813 -3580 -3789 -3556
rect -3572 -3563 -3547 -3540
rect -3529 -3563 -3504 -3542
rect -3487 -3563 -3462 -3540
rect -3431 -3560 -3374 -3535
rect -3356 -3563 -3331 -3540
rect -3313 -3563 -3288 -3542
rect -3271 -3563 -3246 -3540
rect -3215 -3560 -3158 -3535
rect -6090 -3642 -6066 -3618
rect -6051 -3628 -6017 -3622
rect -6051 -3658 -5989 -3628
rect -4299 -3657 -4275 -3605
rect -3809 -3653 -3785 -3629
rect -3770 -3639 -3736 -3633
rect -6023 -3664 -5989 -3658
rect -3770 -3669 -3708 -3639
rect -6090 -3697 -6066 -3673
rect -3742 -3675 -3708 -3669
rect -3809 -3708 -3785 -3684
rect -3585 -3693 -3560 -3670
rect -3542 -3693 -3517 -3672
rect -3500 -3693 -3475 -3670
rect -3444 -3690 -3387 -3665
rect -3369 -3693 -3344 -3670
rect -3326 -3693 -3301 -3672
rect -3284 -3693 -3259 -3670
rect -3228 -3690 -3171 -3665
rect -6087 -3786 -6063 -3762
rect -6048 -3772 -6014 -3766
rect -6048 -3802 -5986 -3772
rect -4300 -3800 -4276 -3748
rect -3808 -3796 -3784 -3772
rect -3769 -3782 -3735 -3776
rect -6020 -3808 -5986 -3802
rect -3769 -3812 -3707 -3782
rect -6087 -3841 -6063 -3817
rect -3741 -3818 -3707 -3812
rect -3808 -3851 -3784 -3827
rect -3584 -3836 -3559 -3813
rect -3541 -3836 -3516 -3815
rect -3499 -3836 -3474 -3813
rect -3443 -3833 -3386 -3808
rect -3368 -3836 -3343 -3813
rect -3325 -3836 -3300 -3815
rect -3283 -3836 -3258 -3813
rect -3227 -3833 -3170 -3808
rect -6091 -3934 -6067 -3910
rect -6052 -3920 -6018 -3914
rect -6052 -3950 -5990 -3920
rect -6024 -3956 -5990 -3950
rect -4300 -3952 -4276 -3900
rect -3599 -3954 -3574 -3931
rect -3556 -3954 -3531 -3933
rect -3514 -3954 -3489 -3931
rect -3458 -3951 -3401 -3926
rect -3383 -3954 -3358 -3931
rect -3340 -3954 -3315 -3933
rect -3298 -3954 -3273 -3931
rect -3242 -3951 -3185 -3926
rect -6091 -3989 -6067 -3965
rect -6066 -4150 -6042 -4126
rect -6027 -4136 -5993 -4130
rect -6027 -4166 -5965 -4136
rect -5999 -4172 -5965 -4166
rect -6066 -4205 -6042 -4181
rect -6067 -4401 -6031 -4361
rect -6025 -4408 -6001 -4368
rect -6066 -4510 -6030 -4470
rect -6024 -4517 -6000 -4477
rect -6063 -4638 -6027 -4598
rect -6021 -4645 -5997 -4605
rect -6061 -4758 -6025 -4718
rect -6019 -4765 -5995 -4725
rect -6059 -4899 -6023 -4859
rect -6017 -4906 -5993 -4866
rect -5237 -4918 -5213 -4866
<< ntransistor >>
rect -7711 -2630 -7707 -2628
rect -8129 -2636 -8125 -2634
rect -6974 -2632 -6970 -2630
rect -7845 -2637 -7841 -2635
rect -7576 -2636 -7572 -2634
rect -7456 -2635 -7452 -2633
rect -7336 -2635 -7332 -2633
rect -7211 -2634 -7207 -2632
rect -7093 -2634 -7089 -2632
rect -7987 -2639 -7983 -2637
rect -7712 -2673 -7708 -2671
rect -8130 -2679 -8126 -2677
rect -7846 -2680 -7842 -2678
rect -7577 -2679 -7573 -2677
rect -7457 -2678 -7453 -2676
rect -7337 -2678 -7333 -2676
rect -7212 -2677 -7208 -2675
rect -6975 -2675 -6971 -2673
rect -7094 -2677 -7090 -2675
rect -7988 -2682 -7984 -2680
rect -7711 -2715 -7707 -2713
rect -8129 -2721 -8125 -2719
rect -6974 -2717 -6970 -2715
rect -7845 -2722 -7841 -2720
rect -7576 -2721 -7572 -2719
rect -7456 -2720 -7452 -2718
rect -7336 -2720 -7332 -2718
rect -7211 -2719 -7207 -2717
rect -7093 -2719 -7089 -2717
rect -7987 -2724 -7983 -2722
rect -7714 -2776 -7710 -2774
rect -8132 -2782 -8128 -2780
rect -6977 -2778 -6973 -2776
rect -7848 -2783 -7844 -2781
rect -7579 -2782 -7575 -2780
rect -7459 -2781 -7455 -2779
rect -7339 -2781 -7335 -2779
rect -7214 -2780 -7210 -2778
rect -7096 -2780 -7092 -2778
rect -7990 -2785 -7986 -2783
rect -7714 -2797 -7710 -2795
rect -8132 -2803 -8128 -2801
rect -7848 -2804 -7844 -2802
rect -7579 -2803 -7575 -2801
rect -7459 -2802 -7455 -2800
rect -7339 -2802 -7335 -2800
rect -7214 -2801 -7210 -2799
rect -6977 -2799 -6973 -2797
rect -7096 -2801 -7092 -2799
rect -7990 -2806 -7986 -2804
rect -7711 -2846 -7707 -2844
rect -8129 -2852 -8125 -2850
rect -6974 -2848 -6970 -2846
rect -7845 -2853 -7841 -2851
rect -7576 -2852 -7572 -2850
rect -7456 -2851 -7452 -2849
rect -7336 -2851 -7332 -2849
rect -7211 -2850 -7207 -2848
rect -7093 -2850 -7089 -2848
rect -7987 -2855 -7983 -2853
rect -7712 -2889 -7708 -2887
rect -8130 -2895 -8126 -2893
rect -7846 -2896 -7842 -2894
rect -7577 -2895 -7573 -2893
rect -7457 -2894 -7453 -2892
rect -7337 -2894 -7333 -2892
rect -7212 -2893 -7208 -2891
rect -6975 -2891 -6971 -2889
rect -7094 -2893 -7090 -2891
rect -7988 -2898 -7984 -2896
rect -7711 -2931 -7707 -2929
rect -8129 -2937 -8125 -2935
rect -6974 -2933 -6970 -2931
rect -7845 -2938 -7841 -2936
rect -7576 -2937 -7572 -2935
rect -7456 -2936 -7452 -2934
rect -7336 -2936 -7332 -2934
rect -7211 -2935 -7207 -2933
rect -7093 -2935 -7089 -2933
rect -7987 -2940 -7983 -2938
rect -7714 -2992 -7710 -2990
rect -8132 -2998 -8128 -2996
rect -6977 -2994 -6973 -2992
rect -7848 -2999 -7844 -2997
rect -7579 -2998 -7575 -2996
rect -7459 -2997 -7455 -2995
rect -7339 -2997 -7335 -2995
rect -7214 -2996 -7210 -2994
rect -7096 -2996 -7092 -2994
rect -7990 -3001 -7986 -2999
rect -7714 -3013 -7710 -3011
rect -8132 -3019 -8128 -3017
rect -7848 -3020 -7844 -3018
rect -7579 -3019 -7575 -3017
rect -7459 -3018 -7455 -3016
rect -7339 -3018 -7335 -3016
rect -7214 -3017 -7210 -3015
rect -6977 -3015 -6973 -3013
rect -7096 -3017 -7092 -3015
rect -7990 -3022 -7986 -3020
rect -5232 -3068 -5230 -3048
rect -3728 -3225 -3726 -3219
rect -3553 -3260 -3551 -3256
rect -3689 -3274 -3687 -3262
rect -3679 -3274 -3677 -3262
rect -3661 -3274 -3659 -3262
rect -3651 -3274 -3649 -3262
rect -3510 -3261 -3508 -3257
rect -3468 -3260 -3466 -3256
rect -3728 -3280 -3726 -3274
rect -3407 -3263 -3405 -3259
rect -3386 -3263 -3384 -3259
rect -3337 -3260 -3335 -3256
rect -3294 -3261 -3292 -3257
rect -3252 -3260 -3250 -3256
rect -3191 -3263 -3189 -3259
rect -3170 -3263 -3168 -3259
rect -6072 -3484 -6070 -3478
rect -5090 -3499 -5088 -3399
rect -4289 -3427 -4287 -3407
rect -3797 -3409 -3795 -3403
rect -3558 -3444 -3556 -3440
rect -3758 -3458 -3756 -3446
rect -3748 -3458 -3746 -3446
rect -3730 -3458 -3728 -3446
rect -3720 -3458 -3718 -3446
rect -3515 -3445 -3513 -3441
rect -3473 -3444 -3471 -3440
rect -3797 -3464 -3795 -3458
rect -3412 -3447 -3410 -3443
rect -3391 -3447 -3389 -3443
rect -3342 -3444 -3340 -3440
rect -3299 -3445 -3297 -3441
rect -3257 -3444 -3255 -3440
rect -3196 -3447 -3194 -3443
rect -3175 -3447 -3173 -3443
rect -6033 -3533 -6031 -3521
rect -6023 -3533 -6021 -3521
rect -6005 -3533 -6003 -3521
rect -5995 -3533 -5993 -3521
rect -6072 -3539 -6070 -3533
rect -4918 -3588 -4916 -3488
rect -4288 -3558 -4286 -3538
rect -3802 -3539 -3800 -3533
rect -3561 -3575 -3559 -3571
rect -3763 -3588 -3761 -3576
rect -3753 -3588 -3751 -3576
rect -3735 -3588 -3733 -3576
rect -3725 -3588 -3723 -3576
rect -3518 -3576 -3516 -3572
rect -3476 -3575 -3474 -3571
rect -3802 -3594 -3800 -3588
rect -3415 -3578 -3413 -3574
rect -3394 -3578 -3392 -3574
rect -3345 -3575 -3343 -3571
rect -3302 -3576 -3300 -3572
rect -3260 -3575 -3258 -3571
rect -3199 -3578 -3197 -3574
rect -3178 -3578 -3176 -3574
rect -6079 -3656 -6077 -3650
rect -6040 -3705 -6038 -3693
rect -6030 -3705 -6028 -3693
rect -6012 -3705 -6010 -3693
rect -6002 -3705 -6000 -3693
rect -6079 -3711 -6077 -3705
rect -5082 -3767 -5080 -3667
rect -3798 -3667 -3796 -3661
rect -4288 -3689 -4286 -3669
rect -3759 -3716 -3757 -3704
rect -3749 -3716 -3747 -3704
rect -3731 -3716 -3729 -3704
rect -3721 -3716 -3719 -3704
rect -3574 -3705 -3572 -3701
rect -3531 -3706 -3529 -3702
rect -3489 -3705 -3487 -3701
rect -3798 -3722 -3796 -3716
rect -3428 -3708 -3426 -3704
rect -3407 -3708 -3405 -3704
rect -3358 -3705 -3356 -3701
rect -3315 -3706 -3313 -3702
rect -3273 -3705 -3271 -3701
rect -6076 -3800 -6074 -3794
rect -4744 -3822 -4742 -3722
rect -3212 -3708 -3210 -3704
rect -3191 -3708 -3189 -3704
rect -6037 -3849 -6035 -3837
rect -6027 -3849 -6025 -3837
rect -6009 -3849 -6007 -3837
rect -5999 -3849 -5997 -3837
rect -6076 -3855 -6074 -3849
rect -4620 -3853 -4618 -3753
rect -3797 -3810 -3795 -3804
rect -4289 -3832 -4287 -3812
rect -3758 -3859 -3756 -3847
rect -3748 -3859 -3746 -3847
rect -3730 -3859 -3728 -3847
rect -3720 -3859 -3718 -3847
rect -3573 -3848 -3571 -3844
rect -3530 -3849 -3528 -3845
rect -3488 -3848 -3486 -3844
rect -3797 -3865 -3795 -3859
rect -3427 -3851 -3425 -3847
rect -3406 -3851 -3404 -3847
rect -3357 -3848 -3355 -3844
rect -3314 -3849 -3312 -3845
rect -3272 -3848 -3270 -3844
rect -3211 -3851 -3209 -3847
rect -3190 -3851 -3188 -3847
rect -6080 -3948 -6078 -3942
rect -6041 -3997 -6039 -3985
rect -6031 -3997 -6029 -3985
rect -6013 -3997 -6011 -3985
rect -6003 -3997 -6001 -3985
rect -6080 -4003 -6078 -3997
rect -4480 -4016 -4478 -3916
rect -4289 -3984 -4287 -3964
rect -3588 -3966 -3586 -3962
rect -3545 -3967 -3543 -3963
rect -3503 -3966 -3501 -3962
rect -3442 -3969 -3440 -3965
rect -3421 -3969 -3419 -3965
rect -3372 -3966 -3370 -3962
rect -3329 -3967 -3327 -3963
rect -3287 -3966 -3285 -3962
rect -3226 -3969 -3224 -3965
rect -3205 -3969 -3203 -3965
rect -6055 -4164 -6053 -4158
rect -6016 -4213 -6014 -4201
rect -6006 -4213 -6004 -4201
rect -5988 -4213 -5986 -4201
rect -5978 -4213 -5976 -4201
rect -6055 -4219 -6053 -4213
rect -4909 -4391 -4907 -4291
rect -6056 -4444 -6054 -4424
rect -6045 -4444 -6043 -4424
rect -6014 -4426 -6012 -4416
rect -4735 -4424 -4733 -4324
rect -4611 -4495 -4609 -4395
rect -6055 -4553 -6053 -4533
rect -6044 -4553 -6042 -4533
rect -6013 -4535 -6011 -4525
rect -4472 -4594 -4470 -4494
rect -4393 -4653 -4391 -4553
rect -6052 -4681 -6050 -4661
rect -6041 -4681 -6039 -4661
rect -6010 -4663 -6008 -4653
rect -6050 -4801 -6048 -4781
rect -6039 -4801 -6037 -4781
rect -6008 -4783 -6006 -4773
rect -5073 -4911 -5071 -4811
rect -6048 -4942 -6046 -4922
rect -6037 -4942 -6035 -4922
rect -6006 -4924 -6004 -4914
rect -5226 -4950 -5224 -4930
<< ptransistor >>
rect -7692 -2630 -7684 -2628
rect -8110 -2636 -8102 -2634
rect -6955 -2632 -6947 -2630
rect -7826 -2637 -7818 -2635
rect -7557 -2636 -7549 -2634
rect -7437 -2635 -7429 -2633
rect -7317 -2635 -7309 -2633
rect -7192 -2634 -7184 -2632
rect -7074 -2634 -7066 -2632
rect -7968 -2639 -7960 -2637
rect -7692 -2673 -7684 -2671
rect -8110 -2679 -8102 -2677
rect -7826 -2680 -7818 -2678
rect -7557 -2679 -7549 -2677
rect -7437 -2678 -7429 -2676
rect -7317 -2678 -7309 -2676
rect -7192 -2677 -7184 -2675
rect -6955 -2675 -6947 -2673
rect -7074 -2677 -7066 -2675
rect -7968 -2682 -7960 -2680
rect -7692 -2715 -7684 -2713
rect -8110 -2721 -8102 -2719
rect -6955 -2717 -6947 -2715
rect -7826 -2722 -7818 -2720
rect -7557 -2721 -7549 -2719
rect -7437 -2720 -7429 -2718
rect -7317 -2720 -7309 -2718
rect -7192 -2719 -7184 -2717
rect -7074 -2719 -7066 -2717
rect -7968 -2724 -7960 -2722
rect -7689 -2776 -7681 -2774
rect -8107 -2782 -8099 -2780
rect -6952 -2778 -6944 -2776
rect -7823 -2783 -7815 -2781
rect -7554 -2782 -7546 -2780
rect -7434 -2781 -7426 -2779
rect -7314 -2781 -7306 -2779
rect -7189 -2780 -7181 -2778
rect -7071 -2780 -7063 -2778
rect -7965 -2785 -7957 -2783
rect -7689 -2797 -7681 -2795
rect -8107 -2803 -8099 -2801
rect -7823 -2804 -7815 -2802
rect -7554 -2803 -7546 -2801
rect -7434 -2802 -7426 -2800
rect -7314 -2802 -7306 -2800
rect -7189 -2801 -7181 -2799
rect -6952 -2799 -6944 -2797
rect -7071 -2801 -7063 -2799
rect -7965 -2806 -7957 -2804
rect -7692 -2846 -7684 -2844
rect -8110 -2852 -8102 -2850
rect -6955 -2848 -6947 -2846
rect -7826 -2853 -7818 -2851
rect -7557 -2852 -7549 -2850
rect -7437 -2851 -7429 -2849
rect -7317 -2851 -7309 -2849
rect -7192 -2850 -7184 -2848
rect -7074 -2850 -7066 -2848
rect -7968 -2855 -7960 -2853
rect -7692 -2889 -7684 -2887
rect -8110 -2895 -8102 -2893
rect -7826 -2896 -7818 -2894
rect -7557 -2895 -7549 -2893
rect -7437 -2894 -7429 -2892
rect -7317 -2894 -7309 -2892
rect -7192 -2893 -7184 -2891
rect -6955 -2891 -6947 -2889
rect -7074 -2893 -7066 -2891
rect -7968 -2898 -7960 -2896
rect -7692 -2931 -7684 -2929
rect -8110 -2937 -8102 -2935
rect -6955 -2933 -6947 -2931
rect -7826 -2938 -7818 -2936
rect -7557 -2937 -7549 -2935
rect -7437 -2936 -7429 -2934
rect -7317 -2936 -7309 -2934
rect -7192 -2935 -7184 -2933
rect -7074 -2935 -7066 -2933
rect -7968 -2940 -7960 -2938
rect -7689 -2992 -7681 -2990
rect -8107 -2998 -8099 -2996
rect -6952 -2994 -6944 -2992
rect -7823 -2999 -7815 -2997
rect -7554 -2998 -7546 -2996
rect -7434 -2997 -7426 -2995
rect -7314 -2997 -7306 -2995
rect -7189 -2996 -7181 -2994
rect -7071 -2996 -7063 -2994
rect -7965 -3001 -7957 -2999
rect -7689 -3013 -7681 -3011
rect -8107 -3019 -8099 -3017
rect -7823 -3020 -7815 -3018
rect -7554 -3019 -7546 -3017
rect -7434 -3018 -7426 -3016
rect -7314 -3018 -7306 -3016
rect -7189 -3017 -7181 -3015
rect -6952 -3015 -6944 -3013
rect -7071 -3017 -7063 -3015
rect -7965 -3022 -7957 -3020
rect -5232 -3030 -5230 -2990
rect -3728 -3205 -3726 -3193
rect -5098 -3267 -5096 -3217
rect -4926 -3268 -4924 -3218
rect -4752 -3268 -4750 -3218
rect -4628 -3269 -4626 -3219
rect -4488 -3272 -4486 -3222
rect -3689 -3221 -3687 -3197
rect -3679 -3221 -3677 -3197
rect -3661 -3227 -3659 -3203
rect -3651 -3227 -3649 -3203
rect -3728 -3260 -3726 -3248
rect -3553 -3241 -3551 -3233
rect -3510 -3241 -3508 -3233
rect -3468 -3241 -3466 -3233
rect -3407 -3238 -3405 -3230
rect -3386 -3238 -3384 -3230
rect -3337 -3241 -3335 -3233
rect -3294 -3241 -3292 -3233
rect -3252 -3241 -3250 -3233
rect -3191 -3238 -3189 -3230
rect -3170 -3238 -3168 -3230
rect -4289 -3389 -4287 -3349
rect -3797 -3389 -3795 -3377
rect -6072 -3464 -6070 -3452
rect -6033 -3480 -6031 -3456
rect -6023 -3480 -6021 -3456
rect -6005 -3486 -6003 -3462
rect -5995 -3486 -5993 -3462
rect -6072 -3519 -6070 -3507
rect -3758 -3405 -3756 -3381
rect -3748 -3405 -3746 -3381
rect -3730 -3411 -3728 -3387
rect -3720 -3411 -3718 -3387
rect -3797 -3444 -3795 -3432
rect -3558 -3425 -3556 -3417
rect -3515 -3425 -3513 -3417
rect -3473 -3425 -3471 -3417
rect -3412 -3422 -3410 -3414
rect -3391 -3422 -3389 -3414
rect -3342 -3425 -3340 -3417
rect -3299 -3425 -3297 -3417
rect -3257 -3425 -3255 -3417
rect -3196 -3422 -3194 -3414
rect -3175 -3422 -3173 -3414
rect -4288 -3520 -4286 -3480
rect -3802 -3519 -3800 -3507
rect -3763 -3535 -3761 -3511
rect -3753 -3535 -3751 -3511
rect -3735 -3541 -3733 -3517
rect -3725 -3541 -3723 -3517
rect -3802 -3574 -3800 -3562
rect -3561 -3556 -3559 -3548
rect -3518 -3556 -3516 -3548
rect -3476 -3556 -3474 -3548
rect -3415 -3553 -3413 -3545
rect -3394 -3553 -3392 -3545
rect -3345 -3556 -3343 -3548
rect -3302 -3556 -3300 -3548
rect -3260 -3556 -3258 -3548
rect -3199 -3553 -3197 -3545
rect -3178 -3553 -3176 -3545
rect -6079 -3636 -6077 -3624
rect -6040 -3652 -6038 -3628
rect -6030 -3652 -6028 -3628
rect -6012 -3658 -6010 -3634
rect -6002 -3658 -6000 -3634
rect -4288 -3651 -4286 -3611
rect -3798 -3647 -3796 -3635
rect -6079 -3691 -6077 -3679
rect -3759 -3663 -3757 -3639
rect -3749 -3663 -3747 -3639
rect -3731 -3669 -3729 -3645
rect -3721 -3669 -3719 -3645
rect -3798 -3702 -3796 -3690
rect -3574 -3686 -3572 -3678
rect -3531 -3686 -3529 -3678
rect -3489 -3686 -3487 -3678
rect -3428 -3683 -3426 -3675
rect -3407 -3683 -3405 -3675
rect -3358 -3686 -3356 -3678
rect -3315 -3686 -3313 -3678
rect -3273 -3686 -3271 -3678
rect -3212 -3683 -3210 -3675
rect -3191 -3683 -3189 -3675
rect -6076 -3780 -6074 -3768
rect -6037 -3796 -6035 -3772
rect -6027 -3796 -6025 -3772
rect -6009 -3802 -6007 -3778
rect -5999 -3802 -5997 -3778
rect -6076 -3835 -6074 -3823
rect -4289 -3794 -4287 -3754
rect -3797 -3790 -3795 -3778
rect -3758 -3806 -3756 -3782
rect -3748 -3806 -3746 -3782
rect -3730 -3812 -3728 -3788
rect -3720 -3812 -3718 -3788
rect -3797 -3845 -3795 -3833
rect -3573 -3829 -3571 -3821
rect -3530 -3829 -3528 -3821
rect -3488 -3829 -3486 -3821
rect -3427 -3826 -3425 -3818
rect -3406 -3826 -3404 -3818
rect -3357 -3829 -3355 -3821
rect -3314 -3829 -3312 -3821
rect -3272 -3829 -3270 -3821
rect -3211 -3826 -3209 -3818
rect -3190 -3826 -3188 -3818
rect -6080 -3928 -6078 -3916
rect -6041 -3944 -6039 -3920
rect -6031 -3944 -6029 -3920
rect -6013 -3950 -6011 -3926
rect -6003 -3950 -6001 -3926
rect -6080 -3983 -6078 -3971
rect -4289 -3946 -4287 -3906
rect -3588 -3947 -3586 -3939
rect -3545 -3947 -3543 -3939
rect -3503 -3947 -3501 -3939
rect -3442 -3944 -3440 -3936
rect -3421 -3944 -3419 -3936
rect -3372 -3947 -3370 -3939
rect -3329 -3947 -3327 -3939
rect -3287 -3947 -3285 -3939
rect -3226 -3944 -3224 -3936
rect -3205 -3944 -3203 -3936
rect -6055 -4144 -6053 -4132
rect -6016 -4160 -6014 -4136
rect -6006 -4160 -6004 -4136
rect -5988 -4166 -5986 -4142
rect -5978 -4166 -5976 -4142
rect -6055 -4199 -6053 -4187
rect -6056 -4395 -6054 -4375
rect -6045 -4395 -6043 -4375
rect -6014 -4402 -6012 -4382
rect -6055 -4504 -6053 -4484
rect -6044 -4504 -6042 -4484
rect -6013 -4511 -6011 -4491
rect -6052 -4632 -6050 -4612
rect -6041 -4632 -6039 -4612
rect -6010 -4639 -6008 -4619
rect -6050 -4752 -6048 -4732
rect -6039 -4752 -6037 -4732
rect -6008 -4759 -6006 -4739
rect -6048 -4893 -6046 -4873
rect -6037 -4893 -6035 -4873
rect -6006 -4900 -6004 -4880
rect -5226 -4912 -5224 -4872
<< ndiffusion >>
rect -7711 -2628 -7707 -2627
rect -8129 -2634 -8125 -2633
rect -8129 -2637 -8125 -2636
rect -7987 -2637 -7983 -2636
rect -7845 -2635 -7841 -2634
rect -7711 -2631 -7707 -2630
rect -7576 -2634 -7572 -2633
rect -7456 -2633 -7452 -2632
rect -7336 -2633 -7332 -2632
rect -7211 -2632 -7207 -2631
rect -7093 -2632 -7089 -2631
rect -6974 -2630 -6970 -2629
rect -6974 -2633 -6970 -2632
rect -7211 -2635 -7207 -2634
rect -7456 -2636 -7452 -2635
rect -7576 -2637 -7572 -2636
rect -7845 -2638 -7841 -2637
rect -7987 -2640 -7983 -2639
rect -7336 -2636 -7332 -2635
rect -7093 -2635 -7089 -2634
rect -7712 -2671 -7708 -2670
rect -8130 -2677 -8126 -2676
rect -8130 -2680 -8126 -2679
rect -7988 -2680 -7984 -2679
rect -7846 -2678 -7842 -2677
rect -7712 -2674 -7708 -2673
rect -7577 -2677 -7573 -2676
rect -7457 -2676 -7453 -2675
rect -7337 -2676 -7333 -2675
rect -7212 -2675 -7208 -2674
rect -7094 -2675 -7090 -2674
rect -6975 -2673 -6971 -2672
rect -6975 -2676 -6971 -2675
rect -7212 -2678 -7208 -2677
rect -7457 -2679 -7453 -2678
rect -7577 -2680 -7573 -2679
rect -7846 -2681 -7842 -2680
rect -7988 -2683 -7984 -2682
rect -7337 -2679 -7333 -2678
rect -7094 -2678 -7090 -2677
rect -7711 -2713 -7707 -2712
rect -8129 -2719 -8125 -2718
rect -8129 -2722 -8125 -2721
rect -7987 -2722 -7983 -2721
rect -7845 -2720 -7841 -2719
rect -7711 -2716 -7707 -2715
rect -7576 -2719 -7572 -2718
rect -7456 -2718 -7452 -2717
rect -7336 -2718 -7332 -2717
rect -7211 -2717 -7207 -2716
rect -7093 -2717 -7089 -2716
rect -6974 -2715 -6970 -2714
rect -6974 -2718 -6970 -2717
rect -7211 -2720 -7207 -2719
rect -7456 -2721 -7452 -2720
rect -7576 -2722 -7572 -2721
rect -7845 -2723 -7841 -2722
rect -7987 -2725 -7983 -2724
rect -7336 -2721 -7332 -2720
rect -7093 -2720 -7089 -2719
rect -7714 -2774 -7710 -2773
rect -8132 -2780 -8128 -2779
rect -8132 -2783 -8128 -2782
rect -7990 -2783 -7986 -2782
rect -7848 -2781 -7844 -2780
rect -7714 -2777 -7710 -2776
rect -7579 -2780 -7575 -2779
rect -7459 -2779 -7455 -2778
rect -7339 -2779 -7335 -2778
rect -7214 -2778 -7210 -2777
rect -7096 -2778 -7092 -2777
rect -6977 -2776 -6973 -2775
rect -6977 -2779 -6973 -2778
rect -7214 -2781 -7210 -2780
rect -7459 -2782 -7455 -2781
rect -7579 -2783 -7575 -2782
rect -7848 -2784 -7844 -2783
rect -7990 -2786 -7986 -2785
rect -7339 -2782 -7335 -2781
rect -7096 -2781 -7092 -2780
rect -7714 -2795 -7710 -2794
rect -8132 -2801 -8128 -2800
rect -8132 -2804 -8128 -2803
rect -7990 -2804 -7986 -2803
rect -7848 -2802 -7844 -2801
rect -7714 -2798 -7710 -2797
rect -7579 -2801 -7575 -2800
rect -7459 -2800 -7455 -2799
rect -7339 -2800 -7335 -2799
rect -7214 -2799 -7210 -2798
rect -7096 -2799 -7092 -2798
rect -6977 -2797 -6973 -2796
rect -6977 -2800 -6973 -2799
rect -7214 -2802 -7210 -2801
rect -7459 -2803 -7455 -2802
rect -7579 -2804 -7575 -2803
rect -7848 -2805 -7844 -2804
rect -7990 -2807 -7986 -2806
rect -7339 -2803 -7335 -2802
rect -7096 -2802 -7092 -2801
rect -7711 -2844 -7707 -2843
rect -8129 -2850 -8125 -2849
rect -8129 -2853 -8125 -2852
rect -7987 -2853 -7983 -2852
rect -7845 -2851 -7841 -2850
rect -7711 -2847 -7707 -2846
rect -7576 -2850 -7572 -2849
rect -7456 -2849 -7452 -2848
rect -7336 -2849 -7332 -2848
rect -7211 -2848 -7207 -2847
rect -7093 -2848 -7089 -2847
rect -6974 -2846 -6970 -2845
rect -6974 -2849 -6970 -2848
rect -7211 -2851 -7207 -2850
rect -7456 -2852 -7452 -2851
rect -7576 -2853 -7572 -2852
rect -7845 -2854 -7841 -2853
rect -7987 -2856 -7983 -2855
rect -7336 -2852 -7332 -2851
rect -7093 -2851 -7089 -2850
rect -7712 -2887 -7708 -2886
rect -8130 -2893 -8126 -2892
rect -8130 -2896 -8126 -2895
rect -7988 -2896 -7984 -2895
rect -7846 -2894 -7842 -2893
rect -7712 -2890 -7708 -2889
rect -7577 -2893 -7573 -2892
rect -7457 -2892 -7453 -2891
rect -7337 -2892 -7333 -2891
rect -7212 -2891 -7208 -2890
rect -7094 -2891 -7090 -2890
rect -6975 -2889 -6971 -2888
rect -6975 -2892 -6971 -2891
rect -7212 -2894 -7208 -2893
rect -7457 -2895 -7453 -2894
rect -7577 -2896 -7573 -2895
rect -7846 -2897 -7842 -2896
rect -7988 -2899 -7984 -2898
rect -7337 -2895 -7333 -2894
rect -7094 -2894 -7090 -2893
rect -7711 -2929 -7707 -2928
rect -8129 -2935 -8125 -2934
rect -8129 -2938 -8125 -2937
rect -7987 -2938 -7983 -2937
rect -7845 -2936 -7841 -2935
rect -7711 -2932 -7707 -2931
rect -7576 -2935 -7572 -2934
rect -7456 -2934 -7452 -2933
rect -7336 -2934 -7332 -2933
rect -7211 -2933 -7207 -2932
rect -7093 -2933 -7089 -2932
rect -6974 -2931 -6970 -2930
rect -6974 -2934 -6970 -2933
rect -7211 -2936 -7207 -2935
rect -7456 -2937 -7452 -2936
rect -7576 -2938 -7572 -2937
rect -7845 -2939 -7841 -2938
rect -7987 -2941 -7983 -2940
rect -7336 -2937 -7332 -2936
rect -7093 -2936 -7089 -2935
rect -7714 -2990 -7710 -2989
rect -8132 -2996 -8128 -2995
rect -8132 -2999 -8128 -2998
rect -7990 -2999 -7986 -2998
rect -7848 -2997 -7844 -2996
rect -7714 -2993 -7710 -2992
rect -7579 -2996 -7575 -2995
rect -7459 -2995 -7455 -2994
rect -7339 -2995 -7335 -2994
rect -7214 -2994 -7210 -2993
rect -7096 -2994 -7092 -2993
rect -6977 -2992 -6973 -2991
rect -6977 -2995 -6973 -2994
rect -7214 -2997 -7210 -2996
rect -7459 -2998 -7455 -2997
rect -7579 -2999 -7575 -2998
rect -7848 -3000 -7844 -2999
rect -7990 -3002 -7986 -3001
rect -7339 -2998 -7335 -2997
rect -7096 -2997 -7092 -2996
rect -7714 -3011 -7710 -3010
rect -8132 -3017 -8128 -3016
rect -8132 -3020 -8128 -3019
rect -7990 -3020 -7986 -3019
rect -7848 -3018 -7844 -3017
rect -7714 -3014 -7710 -3013
rect -7579 -3017 -7575 -3016
rect -7459 -3016 -7455 -3015
rect -7339 -3016 -7335 -3015
rect -7214 -3015 -7210 -3014
rect -7096 -3015 -7092 -3014
rect -6977 -3013 -6973 -3012
rect -6977 -3016 -6973 -3015
rect -7214 -3018 -7210 -3017
rect -7459 -3019 -7455 -3018
rect -7579 -3020 -7575 -3019
rect -7848 -3021 -7844 -3020
rect -7990 -3023 -7986 -3022
rect -7339 -3019 -7335 -3018
rect -7096 -3018 -7092 -3017
rect -5233 -3068 -5232 -3048
rect -5230 -3068 -5229 -3048
rect -3729 -3225 -3728 -3219
rect -3726 -3225 -3725 -3219
rect -3554 -3260 -3553 -3256
rect -3551 -3260 -3550 -3256
rect -3690 -3274 -3689 -3262
rect -3687 -3274 -3679 -3262
rect -3677 -3274 -3676 -3262
rect -3662 -3274 -3661 -3262
rect -3659 -3274 -3651 -3262
rect -3649 -3274 -3648 -3262
rect -3511 -3261 -3510 -3257
rect -3508 -3261 -3507 -3257
rect -3469 -3260 -3468 -3256
rect -3466 -3260 -3465 -3256
rect -3729 -3280 -3728 -3274
rect -3726 -3280 -3725 -3274
rect -3408 -3263 -3407 -3259
rect -3405 -3263 -3404 -3259
rect -3387 -3263 -3386 -3259
rect -3384 -3263 -3383 -3259
rect -3338 -3260 -3337 -3256
rect -3335 -3260 -3334 -3256
rect -3295 -3261 -3294 -3257
rect -3292 -3261 -3291 -3257
rect -3253 -3260 -3252 -3256
rect -3250 -3260 -3249 -3256
rect -3192 -3263 -3191 -3259
rect -3189 -3263 -3188 -3259
rect -3171 -3263 -3170 -3259
rect -3168 -3263 -3167 -3259
rect -6073 -3484 -6072 -3478
rect -6070 -3484 -6069 -3478
rect -5091 -3499 -5090 -3399
rect -5088 -3499 -5087 -3399
rect -4290 -3427 -4289 -3407
rect -4287 -3427 -4286 -3407
rect -3798 -3409 -3797 -3403
rect -3795 -3409 -3794 -3403
rect -3559 -3444 -3558 -3440
rect -3556 -3444 -3555 -3440
rect -3759 -3458 -3758 -3446
rect -3756 -3458 -3748 -3446
rect -3746 -3458 -3745 -3446
rect -3731 -3458 -3730 -3446
rect -3728 -3458 -3720 -3446
rect -3718 -3458 -3717 -3446
rect -3516 -3445 -3515 -3441
rect -3513 -3445 -3512 -3441
rect -3474 -3444 -3473 -3440
rect -3471 -3444 -3470 -3440
rect -3798 -3464 -3797 -3458
rect -3795 -3464 -3794 -3458
rect -3413 -3447 -3412 -3443
rect -3410 -3447 -3409 -3443
rect -3392 -3447 -3391 -3443
rect -3389 -3447 -3388 -3443
rect -3343 -3444 -3342 -3440
rect -3340 -3444 -3339 -3440
rect -3300 -3445 -3299 -3441
rect -3297 -3445 -3296 -3441
rect -3258 -3444 -3257 -3440
rect -3255 -3444 -3254 -3440
rect -3197 -3447 -3196 -3443
rect -3194 -3447 -3193 -3443
rect -3176 -3447 -3175 -3443
rect -3173 -3447 -3172 -3443
rect -6034 -3533 -6033 -3521
rect -6031 -3533 -6023 -3521
rect -6021 -3533 -6020 -3521
rect -6006 -3533 -6005 -3521
rect -6003 -3533 -5995 -3521
rect -5993 -3533 -5992 -3521
rect -6073 -3539 -6072 -3533
rect -6070 -3539 -6069 -3533
rect -4919 -3588 -4918 -3488
rect -4916 -3588 -4915 -3488
rect -4289 -3558 -4288 -3538
rect -4286 -3558 -4285 -3538
rect -3803 -3539 -3802 -3533
rect -3800 -3539 -3799 -3533
rect -3562 -3575 -3561 -3571
rect -3559 -3575 -3558 -3571
rect -3764 -3588 -3763 -3576
rect -3761 -3588 -3753 -3576
rect -3751 -3588 -3750 -3576
rect -3736 -3588 -3735 -3576
rect -3733 -3588 -3725 -3576
rect -3723 -3588 -3722 -3576
rect -3519 -3576 -3518 -3572
rect -3516 -3576 -3515 -3572
rect -3477 -3575 -3476 -3571
rect -3474 -3575 -3473 -3571
rect -3803 -3594 -3802 -3588
rect -3800 -3594 -3799 -3588
rect -3416 -3578 -3415 -3574
rect -3413 -3578 -3412 -3574
rect -3395 -3578 -3394 -3574
rect -3392 -3578 -3391 -3574
rect -3346 -3575 -3345 -3571
rect -3343 -3575 -3342 -3571
rect -3303 -3576 -3302 -3572
rect -3300 -3576 -3299 -3572
rect -3261 -3575 -3260 -3571
rect -3258 -3575 -3257 -3571
rect -3200 -3578 -3199 -3574
rect -3197 -3578 -3196 -3574
rect -3179 -3578 -3178 -3574
rect -3176 -3578 -3175 -3574
rect -6080 -3656 -6079 -3650
rect -6077 -3656 -6076 -3650
rect -6041 -3705 -6040 -3693
rect -6038 -3705 -6030 -3693
rect -6028 -3705 -6027 -3693
rect -6013 -3705 -6012 -3693
rect -6010 -3705 -6002 -3693
rect -6000 -3705 -5999 -3693
rect -6080 -3711 -6079 -3705
rect -6077 -3711 -6076 -3705
rect -5083 -3767 -5082 -3667
rect -5080 -3767 -5079 -3667
rect -3799 -3667 -3798 -3661
rect -3796 -3667 -3795 -3661
rect -4289 -3689 -4288 -3669
rect -4286 -3689 -4285 -3669
rect -3760 -3716 -3759 -3704
rect -3757 -3716 -3749 -3704
rect -3747 -3716 -3746 -3704
rect -3732 -3716 -3731 -3704
rect -3729 -3716 -3721 -3704
rect -3719 -3716 -3718 -3704
rect -3575 -3705 -3574 -3701
rect -3572 -3705 -3571 -3701
rect -3532 -3706 -3531 -3702
rect -3529 -3706 -3528 -3702
rect -3490 -3705 -3489 -3701
rect -3487 -3705 -3486 -3701
rect -3799 -3722 -3798 -3716
rect -3796 -3722 -3795 -3716
rect -3429 -3708 -3428 -3704
rect -3426 -3708 -3425 -3704
rect -3408 -3708 -3407 -3704
rect -3405 -3708 -3404 -3704
rect -3359 -3705 -3358 -3701
rect -3356 -3705 -3355 -3701
rect -3316 -3706 -3315 -3702
rect -3313 -3706 -3312 -3702
rect -3274 -3705 -3273 -3701
rect -3271 -3705 -3270 -3701
rect -6077 -3800 -6076 -3794
rect -6074 -3800 -6073 -3794
rect -4745 -3822 -4744 -3722
rect -4742 -3822 -4741 -3722
rect -3213 -3708 -3212 -3704
rect -3210 -3708 -3209 -3704
rect -3192 -3708 -3191 -3704
rect -3189 -3708 -3188 -3704
rect -6038 -3849 -6037 -3837
rect -6035 -3849 -6027 -3837
rect -6025 -3849 -6024 -3837
rect -6010 -3849 -6009 -3837
rect -6007 -3849 -5999 -3837
rect -5997 -3849 -5996 -3837
rect -6077 -3855 -6076 -3849
rect -6074 -3855 -6073 -3849
rect -4621 -3853 -4620 -3753
rect -4618 -3853 -4617 -3753
rect -3798 -3810 -3797 -3804
rect -3795 -3810 -3794 -3804
rect -4290 -3832 -4289 -3812
rect -4287 -3832 -4286 -3812
rect -3759 -3859 -3758 -3847
rect -3756 -3859 -3748 -3847
rect -3746 -3859 -3745 -3847
rect -3731 -3859 -3730 -3847
rect -3728 -3859 -3720 -3847
rect -3718 -3859 -3717 -3847
rect -3574 -3848 -3573 -3844
rect -3571 -3848 -3570 -3844
rect -3531 -3849 -3530 -3845
rect -3528 -3849 -3527 -3845
rect -3489 -3848 -3488 -3844
rect -3486 -3848 -3485 -3844
rect -3798 -3865 -3797 -3859
rect -3795 -3865 -3794 -3859
rect -3428 -3851 -3427 -3847
rect -3425 -3851 -3424 -3847
rect -3407 -3851 -3406 -3847
rect -3404 -3851 -3403 -3847
rect -3358 -3848 -3357 -3844
rect -3355 -3848 -3354 -3844
rect -3315 -3849 -3314 -3845
rect -3312 -3849 -3311 -3845
rect -3273 -3848 -3272 -3844
rect -3270 -3848 -3269 -3844
rect -3212 -3851 -3211 -3847
rect -3209 -3851 -3208 -3847
rect -3191 -3851 -3190 -3847
rect -3188 -3851 -3187 -3847
rect -6081 -3948 -6080 -3942
rect -6078 -3948 -6077 -3942
rect -6042 -3997 -6041 -3985
rect -6039 -3997 -6031 -3985
rect -6029 -3997 -6028 -3985
rect -6014 -3997 -6013 -3985
rect -6011 -3997 -6003 -3985
rect -6001 -3997 -6000 -3985
rect -6081 -4003 -6080 -3997
rect -6078 -4003 -6077 -3997
rect -4481 -4016 -4480 -3916
rect -4478 -4016 -4477 -3916
rect -4290 -3984 -4289 -3964
rect -4287 -3984 -4286 -3964
rect -3589 -3966 -3588 -3962
rect -3586 -3966 -3585 -3962
rect -3546 -3967 -3545 -3963
rect -3543 -3967 -3542 -3963
rect -3504 -3966 -3503 -3962
rect -3501 -3966 -3500 -3962
rect -3443 -3969 -3442 -3965
rect -3440 -3969 -3439 -3965
rect -3422 -3969 -3421 -3965
rect -3419 -3969 -3418 -3965
rect -3373 -3966 -3372 -3962
rect -3370 -3966 -3369 -3962
rect -3330 -3967 -3329 -3963
rect -3327 -3967 -3326 -3963
rect -3288 -3966 -3287 -3962
rect -3285 -3966 -3284 -3962
rect -3227 -3969 -3226 -3965
rect -3224 -3969 -3223 -3965
rect -3206 -3969 -3205 -3965
rect -3203 -3969 -3202 -3965
rect -6056 -4164 -6055 -4158
rect -6053 -4164 -6052 -4158
rect -6017 -4213 -6016 -4201
rect -6014 -4213 -6006 -4201
rect -6004 -4213 -6003 -4201
rect -5989 -4213 -5988 -4201
rect -5986 -4213 -5978 -4201
rect -5976 -4213 -5975 -4201
rect -6056 -4219 -6055 -4213
rect -6053 -4219 -6052 -4213
rect -4910 -4391 -4909 -4291
rect -4907 -4391 -4906 -4291
rect -6057 -4444 -6056 -4424
rect -6054 -4444 -6045 -4424
rect -6043 -4444 -6042 -4424
rect -6015 -4426 -6014 -4416
rect -6012 -4426 -6011 -4416
rect -4736 -4424 -4735 -4324
rect -4733 -4424 -4732 -4324
rect -4612 -4495 -4611 -4395
rect -4609 -4495 -4608 -4395
rect -6056 -4553 -6055 -4533
rect -6053 -4553 -6044 -4533
rect -6042 -4553 -6041 -4533
rect -6014 -4535 -6013 -4525
rect -6011 -4535 -6010 -4525
rect -4473 -4594 -4472 -4494
rect -4470 -4594 -4469 -4494
rect -4394 -4653 -4393 -4553
rect -4391 -4653 -4390 -4553
rect -6053 -4681 -6052 -4661
rect -6050 -4681 -6041 -4661
rect -6039 -4681 -6038 -4661
rect -6011 -4663 -6010 -4653
rect -6008 -4663 -6007 -4653
rect -6051 -4801 -6050 -4781
rect -6048 -4801 -6039 -4781
rect -6037 -4801 -6036 -4781
rect -6009 -4783 -6008 -4773
rect -6006 -4783 -6005 -4773
rect -5074 -4911 -5073 -4811
rect -5071 -4911 -5070 -4811
rect -6049 -4942 -6048 -4922
rect -6046 -4942 -6037 -4922
rect -6035 -4942 -6034 -4922
rect -6007 -4924 -6006 -4914
rect -6004 -4924 -6003 -4914
rect -5227 -4950 -5226 -4930
rect -5224 -4950 -5223 -4930
<< pdiffusion >>
rect -7692 -2628 -7684 -2627
rect -8110 -2634 -8102 -2633
rect -8110 -2637 -8102 -2636
rect -7826 -2635 -7818 -2634
rect -7692 -2631 -7684 -2630
rect -7437 -2633 -7429 -2632
rect -7192 -2632 -7184 -2631
rect -6955 -2630 -6947 -2629
rect -7074 -2632 -7066 -2631
rect -7317 -2633 -7309 -2632
rect -7557 -2634 -7549 -2633
rect -7968 -2637 -7960 -2636
rect -7968 -2640 -7960 -2639
rect -7826 -2638 -7818 -2637
rect -7557 -2637 -7549 -2636
rect -7437 -2636 -7429 -2635
rect -7317 -2636 -7309 -2635
rect -7192 -2635 -7184 -2634
rect -7074 -2635 -7066 -2634
rect -6955 -2633 -6947 -2632
rect -7692 -2671 -7684 -2670
rect -8110 -2677 -8102 -2676
rect -8110 -2680 -8102 -2679
rect -7968 -2680 -7960 -2679
rect -7826 -2678 -7818 -2677
rect -7692 -2674 -7684 -2673
rect -7557 -2677 -7549 -2676
rect -7437 -2676 -7429 -2675
rect -7317 -2676 -7309 -2675
rect -7192 -2675 -7184 -2674
rect -7074 -2675 -7066 -2674
rect -6955 -2673 -6947 -2672
rect -7968 -2683 -7960 -2682
rect -7826 -2681 -7818 -2680
rect -7557 -2680 -7549 -2679
rect -7437 -2679 -7429 -2678
rect -7317 -2679 -7309 -2678
rect -7192 -2678 -7184 -2677
rect -7074 -2678 -7066 -2677
rect -6955 -2676 -6947 -2675
rect -7692 -2713 -7684 -2712
rect -8110 -2719 -8102 -2718
rect -8110 -2722 -8102 -2721
rect -7826 -2720 -7818 -2719
rect -7692 -2716 -7684 -2715
rect -7437 -2718 -7429 -2717
rect -7192 -2717 -7184 -2716
rect -6955 -2715 -6947 -2714
rect -7074 -2717 -7066 -2716
rect -7317 -2718 -7309 -2717
rect -7557 -2719 -7549 -2718
rect -7968 -2722 -7960 -2721
rect -7968 -2725 -7960 -2724
rect -7826 -2723 -7818 -2722
rect -7557 -2722 -7549 -2721
rect -7437 -2721 -7429 -2720
rect -7317 -2721 -7309 -2720
rect -7192 -2720 -7184 -2719
rect -7074 -2720 -7066 -2719
rect -6955 -2718 -6947 -2717
rect -7689 -2774 -7681 -2773
rect -8107 -2780 -8099 -2779
rect -8107 -2783 -8099 -2782
rect -7823 -2781 -7815 -2780
rect -7689 -2777 -7681 -2776
rect -7434 -2779 -7426 -2778
rect -7189 -2778 -7181 -2777
rect -6952 -2776 -6944 -2775
rect -7071 -2778 -7063 -2777
rect -7314 -2779 -7306 -2778
rect -7554 -2780 -7546 -2779
rect -7965 -2783 -7957 -2782
rect -7965 -2786 -7957 -2785
rect -7823 -2784 -7815 -2783
rect -7554 -2783 -7546 -2782
rect -7434 -2782 -7426 -2781
rect -7314 -2782 -7306 -2781
rect -7189 -2781 -7181 -2780
rect -7071 -2781 -7063 -2780
rect -6952 -2779 -6944 -2778
rect -7689 -2795 -7681 -2794
rect -8107 -2801 -8099 -2800
rect -8107 -2804 -8099 -2803
rect -7965 -2804 -7957 -2803
rect -7823 -2802 -7815 -2801
rect -7689 -2798 -7681 -2797
rect -7554 -2801 -7546 -2800
rect -7434 -2800 -7426 -2799
rect -7314 -2800 -7306 -2799
rect -7189 -2799 -7181 -2798
rect -7071 -2799 -7063 -2798
rect -6952 -2797 -6944 -2796
rect -7965 -2807 -7957 -2806
rect -7823 -2805 -7815 -2804
rect -7554 -2804 -7546 -2803
rect -7434 -2803 -7426 -2802
rect -7314 -2803 -7306 -2802
rect -7189 -2802 -7181 -2801
rect -7071 -2802 -7063 -2801
rect -6952 -2800 -6944 -2799
rect -7692 -2844 -7684 -2843
rect -8110 -2850 -8102 -2849
rect -8110 -2853 -8102 -2852
rect -7826 -2851 -7818 -2850
rect -7692 -2847 -7684 -2846
rect -7437 -2849 -7429 -2848
rect -7192 -2848 -7184 -2847
rect -6955 -2846 -6947 -2845
rect -7074 -2848 -7066 -2847
rect -7317 -2849 -7309 -2848
rect -7557 -2850 -7549 -2849
rect -7968 -2853 -7960 -2852
rect -7968 -2856 -7960 -2855
rect -7826 -2854 -7818 -2853
rect -7557 -2853 -7549 -2852
rect -7437 -2852 -7429 -2851
rect -7317 -2852 -7309 -2851
rect -7192 -2851 -7184 -2850
rect -7074 -2851 -7066 -2850
rect -6955 -2849 -6947 -2848
rect -7692 -2887 -7684 -2886
rect -8110 -2893 -8102 -2892
rect -8110 -2896 -8102 -2895
rect -7968 -2896 -7960 -2895
rect -7826 -2894 -7818 -2893
rect -7692 -2890 -7684 -2889
rect -7557 -2893 -7549 -2892
rect -7437 -2892 -7429 -2891
rect -7317 -2892 -7309 -2891
rect -7192 -2891 -7184 -2890
rect -7074 -2891 -7066 -2890
rect -6955 -2889 -6947 -2888
rect -7968 -2899 -7960 -2898
rect -7826 -2897 -7818 -2896
rect -7557 -2896 -7549 -2895
rect -7437 -2895 -7429 -2894
rect -7317 -2895 -7309 -2894
rect -7192 -2894 -7184 -2893
rect -7074 -2894 -7066 -2893
rect -6955 -2892 -6947 -2891
rect -7692 -2929 -7684 -2928
rect -8110 -2935 -8102 -2934
rect -8110 -2938 -8102 -2937
rect -7826 -2936 -7818 -2935
rect -7692 -2932 -7684 -2931
rect -7437 -2934 -7429 -2933
rect -7192 -2933 -7184 -2932
rect -6955 -2931 -6947 -2930
rect -7074 -2933 -7066 -2932
rect -7317 -2934 -7309 -2933
rect -7557 -2935 -7549 -2934
rect -7968 -2938 -7960 -2937
rect -7968 -2941 -7960 -2940
rect -7826 -2939 -7818 -2938
rect -7557 -2938 -7549 -2937
rect -7437 -2937 -7429 -2936
rect -7317 -2937 -7309 -2936
rect -7192 -2936 -7184 -2935
rect -7074 -2936 -7066 -2935
rect -6955 -2934 -6947 -2933
rect -7689 -2990 -7681 -2989
rect -8107 -2996 -8099 -2995
rect -8107 -2999 -8099 -2998
rect -7823 -2997 -7815 -2996
rect -7689 -2993 -7681 -2992
rect -7434 -2995 -7426 -2994
rect -7189 -2994 -7181 -2993
rect -6952 -2992 -6944 -2991
rect -7071 -2994 -7063 -2993
rect -7314 -2995 -7306 -2994
rect -7554 -2996 -7546 -2995
rect -7965 -2999 -7957 -2998
rect -7965 -3002 -7957 -3001
rect -7823 -3000 -7815 -2999
rect -7554 -2999 -7546 -2998
rect -7434 -2998 -7426 -2997
rect -7314 -2998 -7306 -2997
rect -7189 -2997 -7181 -2996
rect -7071 -2997 -7063 -2996
rect -6952 -2995 -6944 -2994
rect -7689 -3011 -7681 -3010
rect -8107 -3017 -8099 -3016
rect -8107 -3020 -8099 -3019
rect -7965 -3020 -7957 -3019
rect -7823 -3018 -7815 -3017
rect -7689 -3014 -7681 -3013
rect -7554 -3017 -7546 -3016
rect -7434 -3016 -7426 -3015
rect -7314 -3016 -7306 -3015
rect -7189 -3015 -7181 -3014
rect -7071 -3015 -7063 -3014
rect -6952 -3013 -6944 -3012
rect -7965 -3023 -7957 -3022
rect -7823 -3021 -7815 -3020
rect -7554 -3020 -7546 -3019
rect -7434 -3019 -7426 -3018
rect -7314 -3019 -7306 -3018
rect -7189 -3018 -7181 -3017
rect -7071 -3018 -7063 -3017
rect -6952 -3016 -6944 -3015
rect -5233 -3030 -5232 -2990
rect -5230 -3030 -5229 -2990
rect -3729 -3205 -3728 -3193
rect -3726 -3205 -3725 -3193
rect -5099 -3267 -5098 -3217
rect -5096 -3267 -5095 -3217
rect -4927 -3268 -4926 -3218
rect -4924 -3268 -4923 -3218
rect -4753 -3268 -4752 -3218
rect -4750 -3268 -4749 -3218
rect -4629 -3269 -4628 -3219
rect -4626 -3269 -4625 -3219
rect -4489 -3272 -4488 -3222
rect -4486 -3272 -4485 -3222
rect -3690 -3221 -3689 -3197
rect -3687 -3221 -3685 -3197
rect -3681 -3221 -3679 -3197
rect -3677 -3221 -3676 -3197
rect -3662 -3227 -3661 -3203
rect -3659 -3227 -3657 -3203
rect -3653 -3227 -3651 -3203
rect -3649 -3227 -3648 -3203
rect -3729 -3260 -3728 -3248
rect -3726 -3260 -3725 -3248
rect -3554 -3241 -3553 -3233
rect -3551 -3241 -3550 -3233
rect -3511 -3241 -3510 -3233
rect -3508 -3241 -3507 -3233
rect -3469 -3241 -3468 -3233
rect -3466 -3241 -3465 -3233
rect -3408 -3238 -3407 -3230
rect -3405 -3238 -3404 -3230
rect -3387 -3238 -3386 -3230
rect -3384 -3238 -3383 -3230
rect -3338 -3241 -3337 -3233
rect -3335 -3241 -3334 -3233
rect -3295 -3241 -3294 -3233
rect -3292 -3241 -3291 -3233
rect -3253 -3241 -3252 -3233
rect -3250 -3241 -3249 -3233
rect -3192 -3238 -3191 -3230
rect -3189 -3238 -3188 -3230
rect -3171 -3238 -3170 -3230
rect -3168 -3238 -3167 -3230
rect -4290 -3389 -4289 -3349
rect -4287 -3389 -4286 -3349
rect -3798 -3389 -3797 -3377
rect -3795 -3389 -3794 -3377
rect -6073 -3464 -6072 -3452
rect -6070 -3464 -6069 -3452
rect -6034 -3480 -6033 -3456
rect -6031 -3480 -6029 -3456
rect -6025 -3480 -6023 -3456
rect -6021 -3480 -6020 -3456
rect -6006 -3486 -6005 -3462
rect -6003 -3486 -6001 -3462
rect -5997 -3486 -5995 -3462
rect -5993 -3486 -5992 -3462
rect -6073 -3519 -6072 -3507
rect -6070 -3519 -6069 -3507
rect -3759 -3405 -3758 -3381
rect -3756 -3405 -3754 -3381
rect -3750 -3405 -3748 -3381
rect -3746 -3405 -3745 -3381
rect -3731 -3411 -3730 -3387
rect -3728 -3411 -3726 -3387
rect -3722 -3411 -3720 -3387
rect -3718 -3411 -3717 -3387
rect -3798 -3444 -3797 -3432
rect -3795 -3444 -3794 -3432
rect -3559 -3425 -3558 -3417
rect -3556 -3425 -3555 -3417
rect -3516 -3425 -3515 -3417
rect -3513 -3425 -3512 -3417
rect -3474 -3425 -3473 -3417
rect -3471 -3425 -3470 -3417
rect -3413 -3422 -3412 -3414
rect -3410 -3422 -3409 -3414
rect -3392 -3422 -3391 -3414
rect -3389 -3422 -3388 -3414
rect -3343 -3425 -3342 -3417
rect -3340 -3425 -3339 -3417
rect -3300 -3425 -3299 -3417
rect -3297 -3425 -3296 -3417
rect -3258 -3425 -3257 -3417
rect -3255 -3425 -3254 -3417
rect -3197 -3422 -3196 -3414
rect -3194 -3422 -3193 -3414
rect -3176 -3422 -3175 -3414
rect -3173 -3422 -3172 -3414
rect -4289 -3520 -4288 -3480
rect -4286 -3520 -4285 -3480
rect -3803 -3519 -3802 -3507
rect -3800 -3519 -3799 -3507
rect -3764 -3535 -3763 -3511
rect -3761 -3535 -3759 -3511
rect -3755 -3535 -3753 -3511
rect -3751 -3535 -3750 -3511
rect -3736 -3541 -3735 -3517
rect -3733 -3541 -3731 -3517
rect -3727 -3541 -3725 -3517
rect -3723 -3541 -3722 -3517
rect -3803 -3574 -3802 -3562
rect -3800 -3574 -3799 -3562
rect -3562 -3556 -3561 -3548
rect -3559 -3556 -3558 -3548
rect -3519 -3556 -3518 -3548
rect -3516 -3556 -3515 -3548
rect -3477 -3556 -3476 -3548
rect -3474 -3556 -3473 -3548
rect -3416 -3553 -3415 -3545
rect -3413 -3553 -3412 -3545
rect -3395 -3553 -3394 -3545
rect -3392 -3553 -3391 -3545
rect -3346 -3556 -3345 -3548
rect -3343 -3556 -3342 -3548
rect -3303 -3556 -3302 -3548
rect -3300 -3556 -3299 -3548
rect -3261 -3556 -3260 -3548
rect -3258 -3556 -3257 -3548
rect -3200 -3553 -3199 -3545
rect -3197 -3553 -3196 -3545
rect -3179 -3553 -3178 -3545
rect -3176 -3553 -3175 -3545
rect -6080 -3636 -6079 -3624
rect -6077 -3636 -6076 -3624
rect -6041 -3652 -6040 -3628
rect -6038 -3652 -6036 -3628
rect -6032 -3652 -6030 -3628
rect -6028 -3652 -6027 -3628
rect -6013 -3658 -6012 -3634
rect -6010 -3658 -6008 -3634
rect -6004 -3658 -6002 -3634
rect -6000 -3658 -5999 -3634
rect -4289 -3651 -4288 -3611
rect -4286 -3651 -4285 -3611
rect -3799 -3647 -3798 -3635
rect -3796 -3647 -3795 -3635
rect -6080 -3691 -6079 -3679
rect -6077 -3691 -6076 -3679
rect -3760 -3663 -3759 -3639
rect -3757 -3663 -3755 -3639
rect -3751 -3663 -3749 -3639
rect -3747 -3663 -3746 -3639
rect -3732 -3669 -3731 -3645
rect -3729 -3669 -3727 -3645
rect -3723 -3669 -3721 -3645
rect -3719 -3669 -3718 -3645
rect -3799 -3702 -3798 -3690
rect -3796 -3702 -3795 -3690
rect -3575 -3686 -3574 -3678
rect -3572 -3686 -3571 -3678
rect -3532 -3686 -3531 -3678
rect -3529 -3686 -3528 -3678
rect -3490 -3686 -3489 -3678
rect -3487 -3686 -3486 -3678
rect -3429 -3683 -3428 -3675
rect -3426 -3683 -3425 -3675
rect -3408 -3683 -3407 -3675
rect -3405 -3683 -3404 -3675
rect -3359 -3686 -3358 -3678
rect -3356 -3686 -3355 -3678
rect -3316 -3686 -3315 -3678
rect -3313 -3686 -3312 -3678
rect -3274 -3686 -3273 -3678
rect -3271 -3686 -3270 -3678
rect -3213 -3683 -3212 -3675
rect -3210 -3683 -3209 -3675
rect -3192 -3683 -3191 -3675
rect -3189 -3683 -3188 -3675
rect -6077 -3780 -6076 -3768
rect -6074 -3780 -6073 -3768
rect -6038 -3796 -6037 -3772
rect -6035 -3796 -6033 -3772
rect -6029 -3796 -6027 -3772
rect -6025 -3796 -6024 -3772
rect -6010 -3802 -6009 -3778
rect -6007 -3802 -6005 -3778
rect -6001 -3802 -5999 -3778
rect -5997 -3802 -5996 -3778
rect -6077 -3835 -6076 -3823
rect -6074 -3835 -6073 -3823
rect -4290 -3794 -4289 -3754
rect -4287 -3794 -4286 -3754
rect -3798 -3790 -3797 -3778
rect -3795 -3790 -3794 -3778
rect -3759 -3806 -3758 -3782
rect -3756 -3806 -3754 -3782
rect -3750 -3806 -3748 -3782
rect -3746 -3806 -3745 -3782
rect -3731 -3812 -3730 -3788
rect -3728 -3812 -3726 -3788
rect -3722 -3812 -3720 -3788
rect -3718 -3812 -3717 -3788
rect -3798 -3845 -3797 -3833
rect -3795 -3845 -3794 -3833
rect -3574 -3829 -3573 -3821
rect -3571 -3829 -3570 -3821
rect -3531 -3829 -3530 -3821
rect -3528 -3829 -3527 -3821
rect -3489 -3829 -3488 -3821
rect -3486 -3829 -3485 -3821
rect -3428 -3826 -3427 -3818
rect -3425 -3826 -3424 -3818
rect -3407 -3826 -3406 -3818
rect -3404 -3826 -3403 -3818
rect -3358 -3829 -3357 -3821
rect -3355 -3829 -3354 -3821
rect -3315 -3829 -3314 -3821
rect -3312 -3829 -3311 -3821
rect -3273 -3829 -3272 -3821
rect -3270 -3829 -3269 -3821
rect -3212 -3826 -3211 -3818
rect -3209 -3826 -3208 -3818
rect -3191 -3826 -3190 -3818
rect -3188 -3826 -3187 -3818
rect -6081 -3928 -6080 -3916
rect -6078 -3928 -6077 -3916
rect -6042 -3944 -6041 -3920
rect -6039 -3944 -6037 -3920
rect -6033 -3944 -6031 -3920
rect -6029 -3944 -6028 -3920
rect -6014 -3950 -6013 -3926
rect -6011 -3950 -6009 -3926
rect -6005 -3950 -6003 -3926
rect -6001 -3950 -6000 -3926
rect -6081 -3983 -6080 -3971
rect -6078 -3983 -6077 -3971
rect -4290 -3946 -4289 -3906
rect -4287 -3946 -4286 -3906
rect -3589 -3947 -3588 -3939
rect -3586 -3947 -3585 -3939
rect -3546 -3947 -3545 -3939
rect -3543 -3947 -3542 -3939
rect -3504 -3947 -3503 -3939
rect -3501 -3947 -3500 -3939
rect -3443 -3944 -3442 -3936
rect -3440 -3944 -3439 -3936
rect -3422 -3944 -3421 -3936
rect -3419 -3944 -3418 -3936
rect -3373 -3947 -3372 -3939
rect -3370 -3947 -3369 -3939
rect -3330 -3947 -3329 -3939
rect -3327 -3947 -3326 -3939
rect -3288 -3947 -3287 -3939
rect -3285 -3947 -3284 -3939
rect -3227 -3944 -3226 -3936
rect -3224 -3944 -3223 -3936
rect -3206 -3944 -3205 -3936
rect -3203 -3944 -3202 -3936
rect -6056 -4144 -6055 -4132
rect -6053 -4144 -6052 -4132
rect -6017 -4160 -6016 -4136
rect -6014 -4160 -6012 -4136
rect -6008 -4160 -6006 -4136
rect -6004 -4160 -6003 -4136
rect -5989 -4166 -5988 -4142
rect -5986 -4166 -5984 -4142
rect -5980 -4166 -5978 -4142
rect -5976 -4166 -5975 -4142
rect -6056 -4199 -6055 -4187
rect -6053 -4199 -6052 -4187
rect -6057 -4395 -6056 -4375
rect -6054 -4395 -6050 -4375
rect -6046 -4395 -6045 -4375
rect -6043 -4395 -6042 -4375
rect -6015 -4402 -6014 -4382
rect -6012 -4402 -6011 -4382
rect -6056 -4504 -6055 -4484
rect -6053 -4504 -6049 -4484
rect -6045 -4504 -6044 -4484
rect -6042 -4504 -6041 -4484
rect -6014 -4511 -6013 -4491
rect -6011 -4511 -6010 -4491
rect -6053 -4632 -6052 -4612
rect -6050 -4632 -6046 -4612
rect -6042 -4632 -6041 -4612
rect -6039 -4632 -6038 -4612
rect -6011 -4639 -6010 -4619
rect -6008 -4639 -6007 -4619
rect -6051 -4752 -6050 -4732
rect -6048 -4752 -6044 -4732
rect -6040 -4752 -6039 -4732
rect -6037 -4752 -6036 -4732
rect -6009 -4759 -6008 -4739
rect -6006 -4759 -6005 -4739
rect -6049 -4893 -6048 -4873
rect -6046 -4893 -6042 -4873
rect -6038 -4893 -6037 -4873
rect -6035 -4893 -6034 -4873
rect -6007 -4900 -6006 -4880
rect -6004 -4900 -6003 -4880
rect -5227 -4912 -5226 -4872
rect -5224 -4912 -5223 -4872
<< ndcontact >>
rect -7711 -2627 -7707 -2623
rect -8129 -2633 -8125 -2629
rect -7987 -2636 -7983 -2632
rect -8129 -2641 -8125 -2637
rect -7845 -2634 -7841 -2630
rect -7711 -2635 -7707 -2631
rect -7576 -2633 -7572 -2629
rect -7456 -2632 -7452 -2628
rect -7336 -2632 -7332 -2628
rect -7211 -2631 -7207 -2627
rect -7093 -2631 -7089 -2627
rect -6974 -2629 -6970 -2625
rect -7987 -2644 -7983 -2640
rect -7845 -2642 -7841 -2638
rect -7576 -2641 -7572 -2637
rect -7456 -2640 -7452 -2636
rect -7336 -2640 -7332 -2636
rect -7211 -2639 -7207 -2635
rect -7093 -2639 -7089 -2635
rect -6974 -2637 -6970 -2633
rect -7712 -2670 -7708 -2666
rect -8130 -2676 -8126 -2672
rect -8130 -2684 -8126 -2680
rect -7988 -2679 -7984 -2675
rect -7846 -2677 -7842 -2673
rect -7712 -2678 -7708 -2674
rect -7577 -2676 -7573 -2672
rect -7457 -2675 -7453 -2671
rect -7337 -2675 -7333 -2671
rect -7212 -2674 -7208 -2670
rect -7094 -2674 -7090 -2670
rect -6975 -2672 -6971 -2668
rect -7988 -2687 -7984 -2683
rect -7846 -2685 -7842 -2681
rect -7577 -2684 -7573 -2680
rect -7457 -2683 -7453 -2679
rect -7337 -2683 -7333 -2679
rect -7212 -2682 -7208 -2678
rect -7094 -2682 -7090 -2678
rect -6975 -2680 -6971 -2676
rect -7711 -2712 -7707 -2708
rect -8129 -2718 -8125 -2714
rect -7987 -2721 -7983 -2717
rect -8129 -2726 -8125 -2722
rect -7845 -2719 -7841 -2715
rect -7711 -2720 -7707 -2716
rect -7576 -2718 -7572 -2714
rect -7456 -2717 -7452 -2713
rect -7336 -2717 -7332 -2713
rect -7211 -2716 -7207 -2712
rect -7093 -2716 -7089 -2712
rect -6974 -2714 -6970 -2710
rect -7987 -2729 -7983 -2725
rect -7845 -2727 -7841 -2723
rect -7576 -2726 -7572 -2722
rect -7456 -2725 -7452 -2721
rect -7336 -2725 -7332 -2721
rect -7211 -2724 -7207 -2720
rect -7093 -2724 -7089 -2720
rect -6974 -2722 -6970 -2718
rect -7714 -2773 -7710 -2769
rect -8132 -2779 -8128 -2775
rect -7990 -2782 -7986 -2778
rect -8132 -2787 -8128 -2783
rect -7848 -2780 -7844 -2776
rect -7714 -2781 -7710 -2777
rect -7579 -2779 -7575 -2775
rect -7459 -2778 -7455 -2774
rect -7339 -2778 -7335 -2774
rect -7214 -2777 -7210 -2773
rect -7096 -2777 -7092 -2773
rect -6977 -2775 -6973 -2771
rect -7990 -2790 -7986 -2786
rect -7848 -2788 -7844 -2784
rect -7579 -2787 -7575 -2783
rect -7459 -2786 -7455 -2782
rect -7339 -2786 -7335 -2782
rect -7214 -2785 -7210 -2781
rect -7096 -2785 -7092 -2781
rect -6977 -2783 -6973 -2779
rect -7714 -2794 -7710 -2790
rect -8132 -2800 -8128 -2796
rect -8132 -2808 -8128 -2804
rect -7990 -2803 -7986 -2799
rect -7848 -2801 -7844 -2797
rect -7714 -2802 -7710 -2798
rect -7579 -2800 -7575 -2796
rect -7459 -2799 -7455 -2795
rect -7339 -2799 -7335 -2795
rect -7214 -2798 -7210 -2794
rect -7096 -2798 -7092 -2794
rect -6977 -2796 -6973 -2792
rect -7990 -2811 -7986 -2807
rect -7848 -2809 -7844 -2805
rect -7579 -2808 -7575 -2804
rect -7459 -2807 -7455 -2803
rect -7339 -2807 -7335 -2803
rect -7214 -2806 -7210 -2802
rect -7096 -2806 -7092 -2802
rect -6977 -2804 -6973 -2800
rect -7711 -2843 -7707 -2839
rect -8129 -2849 -8125 -2845
rect -7987 -2852 -7983 -2848
rect -8129 -2857 -8125 -2853
rect -7845 -2850 -7841 -2846
rect -7711 -2851 -7707 -2847
rect -7576 -2849 -7572 -2845
rect -7456 -2848 -7452 -2844
rect -7336 -2848 -7332 -2844
rect -7211 -2847 -7207 -2843
rect -7093 -2847 -7089 -2843
rect -6974 -2845 -6970 -2841
rect -7987 -2860 -7983 -2856
rect -7845 -2858 -7841 -2854
rect -7576 -2857 -7572 -2853
rect -7456 -2856 -7452 -2852
rect -7336 -2856 -7332 -2852
rect -7211 -2855 -7207 -2851
rect -7093 -2855 -7089 -2851
rect -6974 -2853 -6970 -2849
rect -7712 -2886 -7708 -2882
rect -8130 -2892 -8126 -2888
rect -8130 -2900 -8126 -2896
rect -7988 -2895 -7984 -2891
rect -7846 -2893 -7842 -2889
rect -7712 -2894 -7708 -2890
rect -7577 -2892 -7573 -2888
rect -7457 -2891 -7453 -2887
rect -7337 -2891 -7333 -2887
rect -7212 -2890 -7208 -2886
rect -7094 -2890 -7090 -2886
rect -6975 -2888 -6971 -2884
rect -7988 -2903 -7984 -2899
rect -7846 -2901 -7842 -2897
rect -7577 -2900 -7573 -2896
rect -7457 -2899 -7453 -2895
rect -7337 -2899 -7333 -2895
rect -7212 -2898 -7208 -2894
rect -7094 -2898 -7090 -2894
rect -6975 -2896 -6971 -2892
rect -7711 -2928 -7707 -2924
rect -8129 -2934 -8125 -2930
rect -7987 -2937 -7983 -2933
rect -8129 -2942 -8125 -2938
rect -7845 -2935 -7841 -2931
rect -7711 -2936 -7707 -2932
rect -7576 -2934 -7572 -2930
rect -7456 -2933 -7452 -2929
rect -7336 -2933 -7332 -2929
rect -7211 -2932 -7207 -2928
rect -7093 -2932 -7089 -2928
rect -6974 -2930 -6970 -2926
rect -7987 -2945 -7983 -2941
rect -7845 -2943 -7841 -2939
rect -7576 -2942 -7572 -2938
rect -7456 -2941 -7452 -2937
rect -7336 -2941 -7332 -2937
rect -7211 -2940 -7207 -2936
rect -7093 -2940 -7089 -2936
rect -6974 -2938 -6970 -2934
rect -7714 -2989 -7710 -2985
rect -8132 -2995 -8128 -2991
rect -7990 -2998 -7986 -2994
rect -8132 -3003 -8128 -2999
rect -7848 -2996 -7844 -2992
rect -7714 -2997 -7710 -2993
rect -7579 -2995 -7575 -2991
rect -7459 -2994 -7455 -2990
rect -7339 -2994 -7335 -2990
rect -7214 -2993 -7210 -2989
rect -7096 -2993 -7092 -2989
rect -6977 -2991 -6973 -2987
rect -7990 -3006 -7986 -3002
rect -7848 -3004 -7844 -3000
rect -7579 -3003 -7575 -2999
rect -7459 -3002 -7455 -2998
rect -7339 -3002 -7335 -2998
rect -7214 -3001 -7210 -2997
rect -7096 -3001 -7092 -2997
rect -6977 -2999 -6973 -2995
rect -7714 -3010 -7710 -3006
rect -8132 -3016 -8128 -3012
rect -8132 -3024 -8128 -3020
rect -7990 -3019 -7986 -3015
rect -7848 -3017 -7844 -3013
rect -7714 -3018 -7710 -3014
rect -7579 -3016 -7575 -3012
rect -7459 -3015 -7455 -3011
rect -7339 -3015 -7335 -3011
rect -7214 -3014 -7210 -3010
rect -7096 -3014 -7092 -3010
rect -6977 -3012 -6973 -3008
rect -7990 -3027 -7986 -3023
rect -7848 -3025 -7844 -3021
rect -7579 -3024 -7575 -3020
rect -7459 -3023 -7455 -3019
rect -7339 -3023 -7335 -3019
rect -7214 -3022 -7210 -3018
rect -7096 -3022 -7092 -3018
rect -6977 -3020 -6973 -3016
rect -5237 -3068 -5233 -3048
rect -5229 -3068 -5225 -3048
rect -3733 -3225 -3729 -3219
rect -3725 -3225 -3721 -3219
rect -3558 -3260 -3554 -3256
rect -3550 -3260 -3546 -3256
rect -3694 -3274 -3690 -3262
rect -3676 -3274 -3672 -3262
rect -3666 -3274 -3662 -3262
rect -3648 -3274 -3644 -3262
rect -3515 -3261 -3511 -3257
rect -3507 -3261 -3503 -3257
rect -3473 -3260 -3469 -3256
rect -3465 -3260 -3461 -3256
rect -3733 -3280 -3729 -3274
rect -3725 -3280 -3721 -3274
rect -3412 -3263 -3408 -3259
rect -3404 -3263 -3400 -3259
rect -3391 -3263 -3387 -3259
rect -3383 -3263 -3379 -3259
rect -3342 -3260 -3338 -3256
rect -3334 -3260 -3330 -3256
rect -3299 -3261 -3295 -3257
rect -3291 -3261 -3287 -3257
rect -3257 -3260 -3253 -3256
rect -3249 -3260 -3245 -3256
rect -3196 -3263 -3192 -3259
rect -3188 -3263 -3184 -3259
rect -3175 -3263 -3171 -3259
rect -3167 -3263 -3163 -3259
rect -6077 -3484 -6073 -3478
rect -6069 -3484 -6065 -3478
rect -5095 -3499 -5091 -3399
rect -5087 -3499 -5083 -3399
rect -4294 -3427 -4290 -3407
rect -4286 -3427 -4282 -3407
rect -3802 -3409 -3798 -3403
rect -3794 -3409 -3790 -3403
rect -3563 -3444 -3559 -3440
rect -3555 -3444 -3551 -3440
rect -3763 -3458 -3759 -3446
rect -3745 -3458 -3741 -3446
rect -3735 -3458 -3731 -3446
rect -3717 -3458 -3713 -3446
rect -3520 -3445 -3516 -3441
rect -3512 -3445 -3508 -3441
rect -3478 -3444 -3474 -3440
rect -3470 -3444 -3466 -3440
rect -3802 -3464 -3798 -3458
rect -3794 -3464 -3790 -3458
rect -3417 -3447 -3413 -3443
rect -3409 -3447 -3405 -3443
rect -3396 -3447 -3392 -3443
rect -3388 -3447 -3384 -3443
rect -3347 -3444 -3343 -3440
rect -3339 -3444 -3335 -3440
rect -3304 -3445 -3300 -3441
rect -3296 -3445 -3292 -3441
rect -3262 -3444 -3258 -3440
rect -3254 -3444 -3250 -3440
rect -3201 -3447 -3197 -3443
rect -3193 -3447 -3189 -3443
rect -3180 -3447 -3176 -3443
rect -3172 -3447 -3168 -3443
rect -6038 -3533 -6034 -3521
rect -6020 -3533 -6016 -3521
rect -6010 -3533 -6006 -3521
rect -5992 -3533 -5988 -3521
rect -6077 -3539 -6073 -3533
rect -6069 -3539 -6065 -3533
rect -4923 -3588 -4919 -3488
rect -4915 -3588 -4911 -3488
rect -4293 -3558 -4289 -3538
rect -4285 -3558 -4281 -3538
rect -3807 -3539 -3803 -3533
rect -3799 -3539 -3795 -3533
rect -3566 -3575 -3562 -3571
rect -3558 -3575 -3554 -3571
rect -3768 -3588 -3764 -3576
rect -3750 -3588 -3746 -3576
rect -3740 -3588 -3736 -3576
rect -3722 -3588 -3718 -3576
rect -3523 -3576 -3519 -3572
rect -3515 -3576 -3511 -3572
rect -3481 -3575 -3477 -3571
rect -3473 -3575 -3469 -3571
rect -3807 -3594 -3803 -3588
rect -3799 -3594 -3795 -3588
rect -3420 -3578 -3416 -3574
rect -3412 -3578 -3408 -3574
rect -3399 -3578 -3395 -3574
rect -3391 -3578 -3387 -3574
rect -3350 -3575 -3346 -3571
rect -3342 -3575 -3338 -3571
rect -3307 -3576 -3303 -3572
rect -3299 -3576 -3295 -3572
rect -3265 -3575 -3261 -3571
rect -3257 -3575 -3253 -3571
rect -3204 -3578 -3200 -3574
rect -3196 -3578 -3192 -3574
rect -3183 -3578 -3179 -3574
rect -3175 -3578 -3171 -3574
rect -6084 -3656 -6080 -3650
rect -6076 -3656 -6072 -3650
rect -6045 -3705 -6041 -3693
rect -6027 -3705 -6023 -3693
rect -6017 -3705 -6013 -3693
rect -5999 -3705 -5995 -3693
rect -6084 -3711 -6080 -3705
rect -6076 -3711 -6072 -3705
rect -5087 -3767 -5083 -3667
rect -5079 -3767 -5075 -3667
rect -3803 -3667 -3799 -3661
rect -3795 -3667 -3791 -3661
rect -4293 -3689 -4289 -3669
rect -4285 -3689 -4281 -3669
rect -3764 -3716 -3760 -3704
rect -3746 -3716 -3742 -3704
rect -3736 -3716 -3732 -3704
rect -3718 -3716 -3714 -3704
rect -3579 -3705 -3575 -3701
rect -3571 -3705 -3567 -3701
rect -3536 -3706 -3532 -3702
rect -3528 -3706 -3524 -3702
rect -3494 -3705 -3490 -3701
rect -3486 -3705 -3482 -3701
rect -3803 -3722 -3799 -3716
rect -3795 -3722 -3791 -3716
rect -3433 -3708 -3429 -3704
rect -3425 -3708 -3421 -3704
rect -3412 -3708 -3408 -3704
rect -3404 -3708 -3400 -3704
rect -3363 -3705 -3359 -3701
rect -3355 -3705 -3351 -3701
rect -3320 -3706 -3316 -3702
rect -3312 -3706 -3308 -3702
rect -3278 -3705 -3274 -3701
rect -3270 -3705 -3266 -3701
rect -6081 -3800 -6077 -3794
rect -6073 -3800 -6069 -3794
rect -4749 -3822 -4745 -3722
rect -4741 -3822 -4737 -3722
rect -3217 -3708 -3213 -3704
rect -3209 -3708 -3205 -3704
rect -3196 -3708 -3192 -3704
rect -3188 -3708 -3184 -3704
rect -6042 -3849 -6038 -3837
rect -6024 -3849 -6020 -3837
rect -6014 -3849 -6010 -3837
rect -5996 -3849 -5992 -3837
rect -6081 -3855 -6077 -3849
rect -6073 -3855 -6069 -3849
rect -4625 -3853 -4621 -3753
rect -4617 -3853 -4613 -3753
rect -3802 -3810 -3798 -3804
rect -3794 -3810 -3790 -3804
rect -4294 -3832 -4290 -3812
rect -4286 -3832 -4282 -3812
rect -3763 -3859 -3759 -3847
rect -3745 -3859 -3741 -3847
rect -3735 -3859 -3731 -3847
rect -3717 -3859 -3713 -3847
rect -3578 -3848 -3574 -3844
rect -3570 -3848 -3566 -3844
rect -3535 -3849 -3531 -3845
rect -3527 -3849 -3523 -3845
rect -3493 -3848 -3489 -3844
rect -3485 -3848 -3481 -3844
rect -3802 -3865 -3798 -3859
rect -3794 -3865 -3790 -3859
rect -3432 -3851 -3428 -3847
rect -3424 -3851 -3420 -3847
rect -3411 -3851 -3407 -3847
rect -3403 -3851 -3399 -3847
rect -3362 -3848 -3358 -3844
rect -3354 -3848 -3350 -3844
rect -3319 -3849 -3315 -3845
rect -3311 -3849 -3307 -3845
rect -3277 -3848 -3273 -3844
rect -3269 -3848 -3265 -3844
rect -3216 -3851 -3212 -3847
rect -3208 -3851 -3204 -3847
rect -3195 -3851 -3191 -3847
rect -3187 -3851 -3183 -3847
rect -6085 -3948 -6081 -3942
rect -6077 -3948 -6073 -3942
rect -6046 -3997 -6042 -3985
rect -6028 -3997 -6024 -3985
rect -6018 -3997 -6014 -3985
rect -6000 -3997 -5996 -3985
rect -6085 -4003 -6081 -3997
rect -6077 -4003 -6073 -3997
rect -4485 -4016 -4481 -3916
rect -4477 -4016 -4473 -3916
rect -4294 -3984 -4290 -3964
rect -4286 -3984 -4282 -3964
rect -3593 -3966 -3589 -3962
rect -3585 -3966 -3581 -3962
rect -3550 -3967 -3546 -3963
rect -3542 -3967 -3538 -3963
rect -3508 -3966 -3504 -3962
rect -3500 -3966 -3496 -3962
rect -3447 -3969 -3443 -3965
rect -3439 -3969 -3435 -3965
rect -3426 -3969 -3422 -3965
rect -3418 -3969 -3414 -3965
rect -3377 -3966 -3373 -3962
rect -3369 -3966 -3365 -3962
rect -3334 -3967 -3330 -3963
rect -3326 -3967 -3322 -3963
rect -3292 -3966 -3288 -3962
rect -3284 -3966 -3280 -3962
rect -3231 -3969 -3227 -3965
rect -3223 -3969 -3219 -3965
rect -3210 -3969 -3206 -3965
rect -3202 -3969 -3198 -3965
rect -6060 -4164 -6056 -4158
rect -6052 -4164 -6048 -4158
rect -6021 -4213 -6017 -4201
rect -6003 -4213 -5999 -4201
rect -5993 -4213 -5989 -4201
rect -5975 -4213 -5971 -4201
rect -6060 -4219 -6056 -4213
rect -6052 -4219 -6048 -4213
rect -4914 -4391 -4910 -4291
rect -4906 -4391 -4902 -4291
rect -6061 -4444 -6057 -4424
rect -6042 -4444 -6038 -4424
rect -6019 -4426 -6015 -4416
rect -6011 -4426 -6007 -4416
rect -4740 -4424 -4736 -4324
rect -4732 -4424 -4728 -4324
rect -4616 -4495 -4612 -4395
rect -4608 -4495 -4604 -4395
rect -6060 -4553 -6056 -4533
rect -6041 -4553 -6037 -4533
rect -6018 -4535 -6014 -4525
rect -6010 -4535 -6006 -4525
rect -4477 -4594 -4473 -4494
rect -4469 -4594 -4465 -4494
rect -4398 -4653 -4394 -4553
rect -4390 -4653 -4386 -4553
rect -6057 -4681 -6053 -4661
rect -6038 -4681 -6034 -4661
rect -6015 -4663 -6011 -4653
rect -6007 -4663 -6003 -4653
rect -6055 -4801 -6051 -4781
rect -6036 -4801 -6032 -4781
rect -6013 -4783 -6009 -4773
rect -6005 -4783 -6001 -4773
rect -5078 -4911 -5074 -4811
rect -5070 -4911 -5066 -4811
rect -6053 -4942 -6049 -4922
rect -6034 -4942 -6030 -4922
rect -6011 -4924 -6007 -4914
rect -6003 -4924 -5999 -4914
rect -5231 -4950 -5227 -4930
rect -5223 -4950 -5219 -4930
<< pdcontact >>
rect -7692 -2627 -7684 -2623
rect -8110 -2633 -8102 -2629
rect -7968 -2636 -7960 -2632
rect -7826 -2634 -7818 -2630
rect -7692 -2635 -7684 -2631
rect -7557 -2633 -7549 -2629
rect -7437 -2632 -7429 -2628
rect -7317 -2632 -7309 -2628
rect -7192 -2631 -7184 -2627
rect -7074 -2631 -7066 -2627
rect -6955 -2629 -6947 -2625
rect -8110 -2641 -8102 -2637
rect -7968 -2644 -7960 -2640
rect -7826 -2642 -7818 -2638
rect -7557 -2641 -7549 -2637
rect -7437 -2640 -7429 -2636
rect -7317 -2640 -7309 -2636
rect -7192 -2639 -7184 -2635
rect -7074 -2639 -7066 -2635
rect -6955 -2637 -6947 -2633
rect -7692 -2670 -7684 -2666
rect -8110 -2676 -8102 -2672
rect -8110 -2684 -8102 -2680
rect -7968 -2679 -7960 -2675
rect -7826 -2677 -7818 -2673
rect -7692 -2678 -7684 -2674
rect -7557 -2676 -7549 -2672
rect -7437 -2675 -7429 -2671
rect -7317 -2675 -7309 -2671
rect -7192 -2674 -7184 -2670
rect -7074 -2674 -7066 -2670
rect -6955 -2672 -6947 -2668
rect -7968 -2687 -7960 -2683
rect -7826 -2685 -7818 -2681
rect -7557 -2684 -7549 -2680
rect -7437 -2683 -7429 -2679
rect -7317 -2683 -7309 -2679
rect -7192 -2682 -7184 -2678
rect -7074 -2682 -7066 -2678
rect -6955 -2680 -6947 -2676
rect -7692 -2712 -7684 -2708
rect -8110 -2718 -8102 -2714
rect -7968 -2721 -7960 -2717
rect -7826 -2719 -7818 -2715
rect -7692 -2720 -7684 -2716
rect -7557 -2718 -7549 -2714
rect -7437 -2717 -7429 -2713
rect -7317 -2717 -7309 -2713
rect -7192 -2716 -7184 -2712
rect -7074 -2716 -7066 -2712
rect -6955 -2714 -6947 -2710
rect -8110 -2726 -8102 -2722
rect -7968 -2729 -7960 -2725
rect -7826 -2727 -7818 -2723
rect -7557 -2726 -7549 -2722
rect -7437 -2725 -7429 -2721
rect -7317 -2725 -7309 -2721
rect -7192 -2724 -7184 -2720
rect -7074 -2724 -7066 -2720
rect -6955 -2722 -6947 -2718
rect -7689 -2773 -7681 -2769
rect -8107 -2779 -8099 -2775
rect -7965 -2782 -7957 -2778
rect -7823 -2780 -7815 -2776
rect -7689 -2781 -7681 -2777
rect -7554 -2779 -7546 -2775
rect -7434 -2778 -7426 -2774
rect -7314 -2778 -7306 -2774
rect -7189 -2777 -7181 -2773
rect -7071 -2777 -7063 -2773
rect -6952 -2775 -6944 -2771
rect -8107 -2787 -8099 -2783
rect -7965 -2790 -7957 -2786
rect -7823 -2788 -7815 -2784
rect -7554 -2787 -7546 -2783
rect -7434 -2786 -7426 -2782
rect -7314 -2786 -7306 -2782
rect -7189 -2785 -7181 -2781
rect -7071 -2785 -7063 -2781
rect -6952 -2783 -6944 -2779
rect -7689 -2794 -7681 -2790
rect -8107 -2800 -8099 -2796
rect -8107 -2808 -8099 -2804
rect -7965 -2803 -7957 -2799
rect -7823 -2801 -7815 -2797
rect -7689 -2802 -7681 -2798
rect -7554 -2800 -7546 -2796
rect -7434 -2799 -7426 -2795
rect -7314 -2799 -7306 -2795
rect -7189 -2798 -7181 -2794
rect -7071 -2798 -7063 -2794
rect -6952 -2796 -6944 -2792
rect -7965 -2811 -7957 -2807
rect -7823 -2809 -7815 -2805
rect -7554 -2808 -7546 -2804
rect -7434 -2807 -7426 -2803
rect -7314 -2807 -7306 -2803
rect -7189 -2806 -7181 -2802
rect -7071 -2806 -7063 -2802
rect -6952 -2804 -6944 -2800
rect -7692 -2843 -7684 -2839
rect -8110 -2849 -8102 -2845
rect -7968 -2852 -7960 -2848
rect -7826 -2850 -7818 -2846
rect -7692 -2851 -7684 -2847
rect -7557 -2849 -7549 -2845
rect -7437 -2848 -7429 -2844
rect -7317 -2848 -7309 -2844
rect -7192 -2847 -7184 -2843
rect -7074 -2847 -7066 -2843
rect -6955 -2845 -6947 -2841
rect -8110 -2857 -8102 -2853
rect -7968 -2860 -7960 -2856
rect -7826 -2858 -7818 -2854
rect -7557 -2857 -7549 -2853
rect -7437 -2856 -7429 -2852
rect -7317 -2856 -7309 -2852
rect -7192 -2855 -7184 -2851
rect -7074 -2855 -7066 -2851
rect -6955 -2853 -6947 -2849
rect -7692 -2886 -7684 -2882
rect -8110 -2892 -8102 -2888
rect -8110 -2900 -8102 -2896
rect -7968 -2895 -7960 -2891
rect -7826 -2893 -7818 -2889
rect -7692 -2894 -7684 -2890
rect -7557 -2892 -7549 -2888
rect -7437 -2891 -7429 -2887
rect -7317 -2891 -7309 -2887
rect -7192 -2890 -7184 -2886
rect -7074 -2890 -7066 -2886
rect -6955 -2888 -6947 -2884
rect -7968 -2903 -7960 -2899
rect -7826 -2901 -7818 -2897
rect -7557 -2900 -7549 -2896
rect -7437 -2899 -7429 -2895
rect -7317 -2899 -7309 -2895
rect -7192 -2898 -7184 -2894
rect -7074 -2898 -7066 -2894
rect -6955 -2896 -6947 -2892
rect -7692 -2928 -7684 -2924
rect -8110 -2934 -8102 -2930
rect -7968 -2937 -7960 -2933
rect -7826 -2935 -7818 -2931
rect -7692 -2936 -7684 -2932
rect -7557 -2934 -7549 -2930
rect -7437 -2933 -7429 -2929
rect -7317 -2933 -7309 -2929
rect -7192 -2932 -7184 -2928
rect -7074 -2932 -7066 -2928
rect -6955 -2930 -6947 -2926
rect -8110 -2942 -8102 -2938
rect -7968 -2945 -7960 -2941
rect -7826 -2943 -7818 -2939
rect -7557 -2942 -7549 -2938
rect -7437 -2941 -7429 -2937
rect -7317 -2941 -7309 -2937
rect -7192 -2940 -7184 -2936
rect -7074 -2940 -7066 -2936
rect -6955 -2938 -6947 -2934
rect -7689 -2989 -7681 -2985
rect -8107 -2995 -8099 -2991
rect -7965 -2998 -7957 -2994
rect -7823 -2996 -7815 -2992
rect -7689 -2997 -7681 -2993
rect -7554 -2995 -7546 -2991
rect -7434 -2994 -7426 -2990
rect -7314 -2994 -7306 -2990
rect -7189 -2993 -7181 -2989
rect -7071 -2993 -7063 -2989
rect -6952 -2991 -6944 -2987
rect -8107 -3003 -8099 -2999
rect -7965 -3006 -7957 -3002
rect -7823 -3004 -7815 -3000
rect -7554 -3003 -7546 -2999
rect -7434 -3002 -7426 -2998
rect -7314 -3002 -7306 -2998
rect -7189 -3001 -7181 -2997
rect -7071 -3001 -7063 -2997
rect -6952 -2999 -6944 -2995
rect -7689 -3010 -7681 -3006
rect -8107 -3016 -8099 -3012
rect -8107 -3024 -8099 -3020
rect -7965 -3019 -7957 -3015
rect -7823 -3017 -7815 -3013
rect -7689 -3018 -7681 -3014
rect -7554 -3016 -7546 -3012
rect -7434 -3015 -7426 -3011
rect -7314 -3015 -7306 -3011
rect -7189 -3014 -7181 -3010
rect -7071 -3014 -7063 -3010
rect -6952 -3012 -6944 -3008
rect -7965 -3027 -7957 -3023
rect -7823 -3025 -7815 -3021
rect -7554 -3024 -7546 -3020
rect -7434 -3023 -7426 -3019
rect -7314 -3023 -7306 -3019
rect -7189 -3022 -7181 -3018
rect -7071 -3022 -7063 -3018
rect -6952 -3020 -6944 -3016
rect -5237 -3030 -5233 -2990
rect -5229 -3030 -5225 -2990
rect -3733 -3205 -3729 -3193
rect -3725 -3205 -3721 -3193
rect -5103 -3267 -5099 -3217
rect -5095 -3267 -5091 -3217
rect -4931 -3268 -4927 -3218
rect -4923 -3268 -4919 -3218
rect -4757 -3268 -4753 -3218
rect -4749 -3268 -4745 -3218
rect -4633 -3269 -4629 -3219
rect -4625 -3269 -4621 -3219
rect -4493 -3272 -4489 -3222
rect -4485 -3272 -4481 -3222
rect -3694 -3221 -3690 -3197
rect -3685 -3221 -3681 -3197
rect -3676 -3221 -3672 -3197
rect -3666 -3227 -3662 -3203
rect -3657 -3227 -3653 -3203
rect -3648 -3227 -3644 -3203
rect -3733 -3260 -3729 -3248
rect -3725 -3260 -3721 -3248
rect -3558 -3241 -3554 -3233
rect -3550 -3241 -3546 -3233
rect -3515 -3241 -3511 -3233
rect -3507 -3241 -3503 -3233
rect -3473 -3241 -3469 -3233
rect -3465 -3241 -3461 -3233
rect -3412 -3238 -3408 -3230
rect -3404 -3238 -3400 -3230
rect -3391 -3238 -3387 -3230
rect -3383 -3238 -3379 -3230
rect -3342 -3241 -3338 -3233
rect -3334 -3241 -3330 -3233
rect -3299 -3241 -3295 -3233
rect -3291 -3241 -3287 -3233
rect -3257 -3241 -3253 -3233
rect -3249 -3241 -3245 -3233
rect -3196 -3238 -3192 -3230
rect -3188 -3238 -3184 -3230
rect -3175 -3238 -3171 -3230
rect -3167 -3238 -3163 -3230
rect -4294 -3389 -4290 -3349
rect -4286 -3389 -4282 -3349
rect -3802 -3389 -3798 -3377
rect -3794 -3389 -3790 -3377
rect -6077 -3464 -6073 -3452
rect -6069 -3464 -6065 -3452
rect -6038 -3480 -6034 -3456
rect -6029 -3480 -6025 -3456
rect -6020 -3480 -6016 -3456
rect -6010 -3486 -6006 -3462
rect -6001 -3486 -5997 -3462
rect -5992 -3486 -5988 -3462
rect -6077 -3519 -6073 -3507
rect -6069 -3519 -6065 -3507
rect -3763 -3405 -3759 -3381
rect -3754 -3405 -3750 -3381
rect -3745 -3405 -3741 -3381
rect -3735 -3411 -3731 -3387
rect -3726 -3411 -3722 -3387
rect -3717 -3411 -3713 -3387
rect -3802 -3444 -3798 -3432
rect -3794 -3444 -3790 -3432
rect -3563 -3425 -3559 -3417
rect -3555 -3425 -3551 -3417
rect -3520 -3425 -3516 -3417
rect -3512 -3425 -3508 -3417
rect -3478 -3425 -3474 -3417
rect -3470 -3425 -3466 -3417
rect -3417 -3422 -3413 -3414
rect -3409 -3422 -3405 -3414
rect -3396 -3422 -3392 -3414
rect -3388 -3422 -3384 -3414
rect -3347 -3425 -3343 -3417
rect -3339 -3425 -3335 -3417
rect -3304 -3425 -3300 -3417
rect -3296 -3425 -3292 -3417
rect -3262 -3425 -3258 -3417
rect -3254 -3425 -3250 -3417
rect -3201 -3422 -3197 -3414
rect -3193 -3422 -3189 -3414
rect -3180 -3422 -3176 -3414
rect -3172 -3422 -3168 -3414
rect -4293 -3520 -4289 -3480
rect -4285 -3520 -4281 -3480
rect -3807 -3519 -3803 -3507
rect -3799 -3519 -3795 -3507
rect -3768 -3535 -3764 -3511
rect -3759 -3535 -3755 -3511
rect -3750 -3535 -3746 -3511
rect -3740 -3541 -3736 -3517
rect -3731 -3541 -3727 -3517
rect -3722 -3541 -3718 -3517
rect -3807 -3574 -3803 -3562
rect -3799 -3574 -3795 -3562
rect -3566 -3556 -3562 -3548
rect -3558 -3556 -3554 -3548
rect -3523 -3556 -3519 -3548
rect -3515 -3556 -3511 -3548
rect -3481 -3556 -3477 -3548
rect -3473 -3556 -3469 -3548
rect -3420 -3553 -3416 -3545
rect -3412 -3553 -3408 -3545
rect -3399 -3553 -3395 -3545
rect -3391 -3553 -3387 -3545
rect -3350 -3556 -3346 -3548
rect -3342 -3556 -3338 -3548
rect -3307 -3556 -3303 -3548
rect -3299 -3556 -3295 -3548
rect -3265 -3556 -3261 -3548
rect -3257 -3556 -3253 -3548
rect -3204 -3553 -3200 -3545
rect -3196 -3553 -3192 -3545
rect -3183 -3553 -3179 -3545
rect -3175 -3553 -3171 -3545
rect -6084 -3636 -6080 -3624
rect -6076 -3636 -6072 -3624
rect -6045 -3652 -6041 -3628
rect -6036 -3652 -6032 -3628
rect -6027 -3652 -6023 -3628
rect -6017 -3658 -6013 -3634
rect -6008 -3658 -6004 -3634
rect -5999 -3658 -5995 -3634
rect -4293 -3651 -4289 -3611
rect -4285 -3651 -4281 -3611
rect -3803 -3647 -3799 -3635
rect -3795 -3647 -3791 -3635
rect -6084 -3691 -6080 -3679
rect -6076 -3691 -6072 -3679
rect -3764 -3663 -3760 -3639
rect -3755 -3663 -3751 -3639
rect -3746 -3663 -3742 -3639
rect -3736 -3669 -3732 -3645
rect -3727 -3669 -3723 -3645
rect -3718 -3669 -3714 -3645
rect -3803 -3702 -3799 -3690
rect -3795 -3702 -3791 -3690
rect -3579 -3686 -3575 -3678
rect -3571 -3686 -3567 -3678
rect -3536 -3686 -3532 -3678
rect -3528 -3686 -3524 -3678
rect -3494 -3686 -3490 -3678
rect -3486 -3686 -3482 -3678
rect -3433 -3683 -3429 -3675
rect -3425 -3683 -3421 -3675
rect -3412 -3683 -3408 -3675
rect -3404 -3683 -3400 -3675
rect -3363 -3686 -3359 -3678
rect -3355 -3686 -3351 -3678
rect -3320 -3686 -3316 -3678
rect -3312 -3686 -3308 -3678
rect -3278 -3686 -3274 -3678
rect -3270 -3686 -3266 -3678
rect -3217 -3683 -3213 -3675
rect -3209 -3683 -3205 -3675
rect -3196 -3683 -3192 -3675
rect -3188 -3683 -3184 -3675
rect -6081 -3780 -6077 -3768
rect -6073 -3780 -6069 -3768
rect -6042 -3796 -6038 -3772
rect -6033 -3796 -6029 -3772
rect -6024 -3796 -6020 -3772
rect -6014 -3802 -6010 -3778
rect -6005 -3802 -6001 -3778
rect -5996 -3802 -5992 -3778
rect -6081 -3835 -6077 -3823
rect -6073 -3835 -6069 -3823
rect -4294 -3794 -4290 -3754
rect -4286 -3794 -4282 -3754
rect -3802 -3790 -3798 -3778
rect -3794 -3790 -3790 -3778
rect -3763 -3806 -3759 -3782
rect -3754 -3806 -3750 -3782
rect -3745 -3806 -3741 -3782
rect -3735 -3812 -3731 -3788
rect -3726 -3812 -3722 -3788
rect -3717 -3812 -3713 -3788
rect -3802 -3845 -3798 -3833
rect -3794 -3845 -3790 -3833
rect -3578 -3829 -3574 -3821
rect -3570 -3829 -3566 -3821
rect -3535 -3829 -3531 -3821
rect -3527 -3829 -3523 -3821
rect -3493 -3829 -3489 -3821
rect -3485 -3829 -3481 -3821
rect -3432 -3826 -3428 -3818
rect -3424 -3826 -3420 -3818
rect -3411 -3826 -3407 -3818
rect -3403 -3826 -3399 -3818
rect -3362 -3829 -3358 -3821
rect -3354 -3829 -3350 -3821
rect -3319 -3829 -3315 -3821
rect -3311 -3829 -3307 -3821
rect -3277 -3829 -3273 -3821
rect -3269 -3829 -3265 -3821
rect -3216 -3826 -3212 -3818
rect -3208 -3826 -3204 -3818
rect -3195 -3826 -3191 -3818
rect -3187 -3826 -3183 -3818
rect -6085 -3928 -6081 -3916
rect -6077 -3928 -6073 -3916
rect -6046 -3944 -6042 -3920
rect -6037 -3944 -6033 -3920
rect -6028 -3944 -6024 -3920
rect -6018 -3950 -6014 -3926
rect -6009 -3950 -6005 -3926
rect -6000 -3950 -5996 -3926
rect -6085 -3983 -6081 -3971
rect -6077 -3983 -6073 -3971
rect -4294 -3946 -4290 -3906
rect -4286 -3946 -4282 -3906
rect -3593 -3947 -3589 -3939
rect -3585 -3947 -3581 -3939
rect -3550 -3947 -3546 -3939
rect -3542 -3947 -3538 -3939
rect -3508 -3947 -3504 -3939
rect -3500 -3947 -3496 -3939
rect -3447 -3944 -3443 -3936
rect -3439 -3944 -3435 -3936
rect -3426 -3944 -3422 -3936
rect -3418 -3944 -3414 -3936
rect -3377 -3947 -3373 -3939
rect -3369 -3947 -3365 -3939
rect -3334 -3947 -3330 -3939
rect -3326 -3947 -3322 -3939
rect -3292 -3947 -3288 -3939
rect -3284 -3947 -3280 -3939
rect -3231 -3944 -3227 -3936
rect -3223 -3944 -3219 -3936
rect -3210 -3944 -3206 -3936
rect -3202 -3944 -3198 -3936
rect -6060 -4144 -6056 -4132
rect -6052 -4144 -6048 -4132
rect -6021 -4160 -6017 -4136
rect -6012 -4160 -6008 -4136
rect -6003 -4160 -5999 -4136
rect -5993 -4166 -5989 -4142
rect -5984 -4166 -5980 -4142
rect -5975 -4166 -5971 -4142
rect -6060 -4199 -6056 -4187
rect -6052 -4199 -6048 -4187
rect -6061 -4395 -6057 -4375
rect -6050 -4395 -6046 -4375
rect -6042 -4395 -6038 -4375
rect -6019 -4402 -6015 -4382
rect -6011 -4402 -6007 -4382
rect -6060 -4504 -6056 -4484
rect -6049 -4504 -6045 -4484
rect -6041 -4504 -6037 -4484
rect -6018 -4511 -6014 -4491
rect -6010 -4511 -6006 -4491
rect -6057 -4632 -6053 -4612
rect -6046 -4632 -6042 -4612
rect -6038 -4632 -6034 -4612
rect -6015 -4639 -6011 -4619
rect -6007 -4639 -6003 -4619
rect -6055 -4752 -6051 -4732
rect -6044 -4752 -6040 -4732
rect -6036 -4752 -6032 -4732
rect -6013 -4759 -6009 -4739
rect -6005 -4759 -6001 -4739
rect -6053 -4893 -6049 -4873
rect -6042 -4893 -6038 -4873
rect -6034 -4893 -6030 -4873
rect -6011 -4900 -6007 -4880
rect -6003 -4900 -5999 -4880
rect -5231 -4912 -5227 -4872
rect -5223 -4912 -5219 -4872
<< psubstratepcontact >>
rect -6005 -4435 -6000 -4431
rect -6004 -4544 -5999 -4540
rect -6001 -4672 -5996 -4668
rect -5999 -4792 -5994 -4788
rect -5997 -4933 -5992 -4929
<< nsubstratencontact >>
rect -5242 -2984 -5238 -2980
rect -5108 -3211 -5104 -3206
rect -4936 -3212 -4932 -3207
rect -4762 -3212 -4758 -3207
rect -4638 -3213 -4634 -3208
rect -4498 -3216 -4494 -3211
rect -4299 -3343 -4295 -3339
rect -4298 -3474 -4294 -3470
rect -4298 -3605 -4294 -3601
rect -4299 -3748 -4295 -3744
rect -4299 -3900 -4295 -3896
rect -6061 -4370 -6057 -4364
rect -6009 -4375 -6005 -4371
rect -6060 -4479 -6056 -4473
rect -6008 -4484 -6004 -4480
rect -6057 -4607 -6053 -4601
rect -6005 -4612 -6001 -4608
rect -6055 -4727 -6051 -4721
rect -6003 -4732 -5999 -4728
rect -6053 -4868 -6049 -4862
rect -5236 -4866 -5232 -4862
rect -6001 -4873 -5997 -4869
<< polysilicon >>
rect -7714 -2630 -7711 -2628
rect -7707 -2630 -7692 -2628
rect -8132 -2636 -8129 -2634
rect -8125 -2636 -8110 -2634
rect -6977 -2632 -6974 -2630
rect -6970 -2632 -6955 -2630
rect -7848 -2637 -7845 -2635
rect -7841 -2637 -7826 -2635
rect -7579 -2636 -7576 -2634
rect -7572 -2636 -7557 -2634
rect -7459 -2635 -7456 -2633
rect -7452 -2635 -7437 -2633
rect -7339 -2635 -7336 -2633
rect -7332 -2635 -7317 -2633
rect -7214 -2634 -7211 -2632
rect -7207 -2634 -7192 -2632
rect -7096 -2634 -7093 -2632
rect -7089 -2634 -7074 -2632
rect -7990 -2639 -7987 -2637
rect -7983 -2639 -7968 -2637
rect -7726 -2673 -7712 -2671
rect -7708 -2673 -7703 -2671
rect -7699 -2673 -7692 -2671
rect -7682 -2673 -7665 -2671
rect -8144 -2679 -8130 -2677
rect -8126 -2679 -8121 -2677
rect -8117 -2679 -8110 -2677
rect -8100 -2679 -8083 -2677
rect -7860 -2680 -7846 -2678
rect -7842 -2680 -7837 -2678
rect -7833 -2680 -7826 -2678
rect -7816 -2680 -7799 -2678
rect -7591 -2679 -7577 -2677
rect -7573 -2679 -7568 -2677
rect -7564 -2679 -7557 -2677
rect -7547 -2679 -7530 -2677
rect -7471 -2678 -7457 -2676
rect -7453 -2678 -7448 -2676
rect -7444 -2678 -7437 -2676
rect -7427 -2678 -7410 -2676
rect -7351 -2678 -7337 -2676
rect -7333 -2678 -7328 -2676
rect -7324 -2678 -7317 -2676
rect -7307 -2678 -7290 -2676
rect -7226 -2677 -7212 -2675
rect -7208 -2677 -7203 -2675
rect -7199 -2677 -7192 -2675
rect -7182 -2677 -7165 -2675
rect -6989 -2675 -6975 -2673
rect -6971 -2675 -6966 -2673
rect -6962 -2675 -6955 -2673
rect -6945 -2675 -6928 -2673
rect -7108 -2677 -7094 -2675
rect -7090 -2677 -7085 -2675
rect -7081 -2677 -7074 -2675
rect -7064 -2677 -7047 -2675
rect -8002 -2682 -7988 -2680
rect -7984 -2682 -7979 -2680
rect -7975 -2682 -7968 -2680
rect -7958 -2682 -7941 -2680
rect -7714 -2715 -7711 -2713
rect -7707 -2715 -7692 -2713
rect -8132 -2721 -8129 -2719
rect -8125 -2721 -8110 -2719
rect -6977 -2717 -6974 -2715
rect -6970 -2717 -6955 -2715
rect -7848 -2722 -7845 -2720
rect -7841 -2722 -7826 -2720
rect -7579 -2721 -7576 -2719
rect -7572 -2721 -7557 -2719
rect -7459 -2720 -7456 -2718
rect -7452 -2720 -7437 -2718
rect -7339 -2720 -7336 -2718
rect -7332 -2720 -7317 -2718
rect -7214 -2719 -7211 -2717
rect -7207 -2719 -7192 -2717
rect -7096 -2719 -7093 -2717
rect -7089 -2719 -7074 -2717
rect -7990 -2724 -7987 -2722
rect -7983 -2724 -7968 -2722
rect -7717 -2776 -7714 -2774
rect -7710 -2776 -7689 -2774
rect -7680 -2776 -7678 -2774
rect -8135 -2782 -8132 -2780
rect -8128 -2782 -8107 -2780
rect -8098 -2782 -8096 -2780
rect -6980 -2778 -6977 -2776
rect -6973 -2778 -6952 -2776
rect -6943 -2778 -6941 -2776
rect -7851 -2783 -7848 -2781
rect -7844 -2783 -7823 -2781
rect -7814 -2783 -7812 -2781
rect -7582 -2782 -7579 -2780
rect -7575 -2782 -7554 -2780
rect -7545 -2782 -7543 -2780
rect -7462 -2781 -7459 -2779
rect -7455 -2781 -7434 -2779
rect -7425 -2781 -7423 -2779
rect -7342 -2781 -7339 -2779
rect -7335 -2781 -7314 -2779
rect -7305 -2781 -7303 -2779
rect -7217 -2780 -7214 -2778
rect -7210 -2780 -7189 -2778
rect -7180 -2780 -7178 -2778
rect -7099 -2780 -7096 -2778
rect -7092 -2780 -7071 -2778
rect -7062 -2780 -7060 -2778
rect -7993 -2785 -7990 -2783
rect -7986 -2785 -7965 -2783
rect -7956 -2785 -7954 -2783
rect -7730 -2797 -7714 -2795
rect -7710 -2797 -7707 -2795
rect -7693 -2797 -7689 -2795
rect -7681 -2797 -7662 -2795
rect -8148 -2803 -8132 -2801
rect -8128 -2803 -8125 -2801
rect -8111 -2803 -8107 -2801
rect -8099 -2803 -8080 -2801
rect -7864 -2804 -7848 -2802
rect -7844 -2804 -7841 -2802
rect -7827 -2804 -7823 -2802
rect -7815 -2804 -7796 -2802
rect -7595 -2803 -7579 -2801
rect -7575 -2803 -7572 -2801
rect -7558 -2803 -7554 -2801
rect -7546 -2803 -7527 -2801
rect -7475 -2802 -7459 -2800
rect -7455 -2802 -7452 -2800
rect -7438 -2802 -7434 -2800
rect -7426 -2802 -7407 -2800
rect -7355 -2802 -7339 -2800
rect -7335 -2802 -7332 -2800
rect -7318 -2802 -7314 -2800
rect -7306 -2802 -7287 -2800
rect -7230 -2801 -7214 -2799
rect -7210 -2801 -7207 -2799
rect -7193 -2801 -7189 -2799
rect -7181 -2801 -7162 -2799
rect -6993 -2799 -6977 -2797
rect -6973 -2799 -6970 -2797
rect -6956 -2799 -6952 -2797
rect -6944 -2799 -6925 -2797
rect -7112 -2801 -7096 -2799
rect -7092 -2801 -7089 -2799
rect -7075 -2801 -7071 -2799
rect -7063 -2801 -7044 -2799
rect -8006 -2806 -7990 -2804
rect -7986 -2806 -7983 -2804
rect -7969 -2806 -7965 -2804
rect -7957 -2806 -7938 -2804
rect -7714 -2846 -7711 -2844
rect -7707 -2846 -7692 -2844
rect -8132 -2852 -8129 -2850
rect -8125 -2852 -8110 -2850
rect -6977 -2848 -6974 -2846
rect -6970 -2848 -6955 -2846
rect -7848 -2853 -7845 -2851
rect -7841 -2853 -7826 -2851
rect -7579 -2852 -7576 -2850
rect -7572 -2852 -7557 -2850
rect -7459 -2851 -7456 -2849
rect -7452 -2851 -7437 -2849
rect -7339 -2851 -7336 -2849
rect -7332 -2851 -7317 -2849
rect -7214 -2850 -7211 -2848
rect -7207 -2850 -7192 -2848
rect -7096 -2850 -7093 -2848
rect -7089 -2850 -7074 -2848
rect -7990 -2855 -7987 -2853
rect -7983 -2855 -7968 -2853
rect -7726 -2889 -7712 -2887
rect -7708 -2889 -7703 -2887
rect -7699 -2889 -7692 -2887
rect -7682 -2889 -7665 -2887
rect -8144 -2895 -8130 -2893
rect -8126 -2895 -8121 -2893
rect -8117 -2895 -8110 -2893
rect -8100 -2895 -8083 -2893
rect -7860 -2896 -7846 -2894
rect -7842 -2896 -7837 -2894
rect -7833 -2896 -7826 -2894
rect -7816 -2896 -7799 -2894
rect -7591 -2895 -7577 -2893
rect -7573 -2895 -7568 -2893
rect -7564 -2895 -7557 -2893
rect -7547 -2895 -7530 -2893
rect -7471 -2894 -7457 -2892
rect -7453 -2894 -7448 -2892
rect -7444 -2894 -7437 -2892
rect -7427 -2894 -7410 -2892
rect -7351 -2894 -7337 -2892
rect -7333 -2894 -7328 -2892
rect -7324 -2894 -7317 -2892
rect -7307 -2894 -7290 -2892
rect -7226 -2893 -7212 -2891
rect -7208 -2893 -7203 -2891
rect -7199 -2893 -7192 -2891
rect -7182 -2893 -7165 -2891
rect -6989 -2891 -6975 -2889
rect -6971 -2891 -6966 -2889
rect -6962 -2891 -6955 -2889
rect -6945 -2891 -6928 -2889
rect -7108 -2893 -7094 -2891
rect -7090 -2893 -7085 -2891
rect -7081 -2893 -7074 -2891
rect -7064 -2893 -7047 -2891
rect -8002 -2898 -7988 -2896
rect -7984 -2898 -7979 -2896
rect -7975 -2898 -7968 -2896
rect -7958 -2898 -7941 -2896
rect -7714 -2931 -7711 -2929
rect -7707 -2931 -7692 -2929
rect -8132 -2937 -8129 -2935
rect -8125 -2937 -8110 -2935
rect -6977 -2933 -6974 -2931
rect -6970 -2933 -6955 -2931
rect -7848 -2938 -7845 -2936
rect -7841 -2938 -7826 -2936
rect -7579 -2937 -7576 -2935
rect -7572 -2937 -7557 -2935
rect -7459 -2936 -7456 -2934
rect -7452 -2936 -7437 -2934
rect -7339 -2936 -7336 -2934
rect -7332 -2936 -7317 -2934
rect -7214 -2935 -7211 -2933
rect -7207 -2935 -7192 -2933
rect -7096 -2935 -7093 -2933
rect -7089 -2935 -7074 -2933
rect -7990 -2940 -7987 -2938
rect -7983 -2940 -7968 -2938
rect -7717 -2992 -7714 -2990
rect -7710 -2992 -7689 -2990
rect -7680 -2992 -7678 -2990
rect -8135 -2998 -8132 -2996
rect -8128 -2998 -8107 -2996
rect -8098 -2998 -8096 -2996
rect -5232 -2990 -5230 -2987
rect -6980 -2994 -6977 -2992
rect -6973 -2994 -6952 -2992
rect -6943 -2994 -6941 -2992
rect -7851 -2999 -7848 -2997
rect -7844 -2999 -7823 -2997
rect -7814 -2999 -7812 -2997
rect -7582 -2998 -7579 -2996
rect -7575 -2998 -7554 -2996
rect -7545 -2998 -7543 -2996
rect -7462 -2997 -7459 -2995
rect -7455 -2997 -7434 -2995
rect -7425 -2997 -7423 -2995
rect -7342 -2997 -7339 -2995
rect -7335 -2997 -7314 -2995
rect -7305 -2997 -7303 -2995
rect -7217 -2996 -7214 -2994
rect -7210 -2996 -7189 -2994
rect -7180 -2996 -7178 -2994
rect -7099 -2996 -7096 -2994
rect -7092 -2996 -7071 -2994
rect -7062 -2996 -7060 -2994
rect -7993 -3001 -7990 -2999
rect -7986 -3001 -7965 -2999
rect -7956 -3001 -7954 -2999
rect -7730 -3013 -7714 -3011
rect -7710 -3013 -7707 -3011
rect -7693 -3013 -7689 -3011
rect -7681 -3013 -7662 -3011
rect -8148 -3019 -8132 -3017
rect -8128 -3019 -8125 -3017
rect -8111 -3019 -8107 -3017
rect -8099 -3019 -8080 -3017
rect -7864 -3020 -7848 -3018
rect -7844 -3020 -7841 -3018
rect -7827 -3020 -7823 -3018
rect -7815 -3020 -7796 -3018
rect -7595 -3019 -7579 -3017
rect -7575 -3019 -7572 -3017
rect -7558 -3019 -7554 -3017
rect -7546 -3019 -7527 -3017
rect -7475 -3018 -7459 -3016
rect -7455 -3018 -7452 -3016
rect -7438 -3018 -7434 -3016
rect -7426 -3018 -7407 -3016
rect -7355 -3018 -7339 -3016
rect -7335 -3018 -7332 -3016
rect -7318 -3018 -7314 -3016
rect -7306 -3018 -7287 -3016
rect -7230 -3017 -7214 -3015
rect -7210 -3017 -7207 -3015
rect -7193 -3017 -7189 -3015
rect -7181 -3017 -7162 -3015
rect -6993 -3015 -6977 -3013
rect -6973 -3015 -6970 -3013
rect -6956 -3015 -6952 -3013
rect -6944 -3015 -6925 -3013
rect -7112 -3017 -7096 -3015
rect -7092 -3017 -7089 -3015
rect -7075 -3017 -7071 -3015
rect -7063 -3017 -7044 -3015
rect -8006 -3022 -7990 -3020
rect -7986 -3022 -7983 -3020
rect -7969 -3022 -7965 -3020
rect -7957 -3022 -7938 -3020
rect -5232 -3048 -5230 -3030
rect -5232 -3072 -5230 -3068
rect -3728 -3193 -3726 -3190
rect -3689 -3197 -3687 -3194
rect -3679 -3197 -3677 -3194
rect -5098 -3217 -5096 -3214
rect -4926 -3218 -4924 -3215
rect -4752 -3218 -4750 -3215
rect -5098 -3290 -5096 -3267
rect -4628 -3219 -4626 -3216
rect -3728 -3219 -3726 -3205
rect -4926 -3291 -4924 -3268
rect -4752 -3291 -4750 -3268
rect -4488 -3222 -4486 -3219
rect -4628 -3292 -4626 -3269
rect -3661 -3203 -3659 -3200
rect -3651 -3203 -3649 -3200
rect -3728 -3228 -3726 -3225
rect -3689 -3230 -3687 -3221
rect -3679 -3231 -3677 -3221
rect -3728 -3248 -3726 -3245
rect -4488 -3295 -4486 -3272
rect -3728 -3274 -3726 -3260
rect -3689 -3262 -3687 -3235
rect -3679 -3262 -3677 -3236
rect -3661 -3238 -3659 -3227
rect -3661 -3262 -3659 -3242
rect -3651 -3249 -3649 -3227
rect -3510 -3231 -3508 -3214
rect -3407 -3229 -3405 -3227
rect -3386 -3230 -3384 -3211
rect -3294 -3231 -3292 -3214
rect -3191 -3229 -3189 -3227
rect -3170 -3230 -3168 -3211
rect -3651 -3262 -3649 -3253
rect -3553 -3256 -3551 -3241
rect -3510 -3248 -3508 -3241
rect -3510 -3257 -3508 -3252
rect -3468 -3256 -3466 -3241
rect -3553 -3263 -3551 -3260
rect -3407 -3259 -3405 -3238
rect -3386 -3242 -3384 -3238
rect -3337 -3256 -3335 -3241
rect -3294 -3248 -3292 -3241
rect -3386 -3259 -3384 -3256
rect -3689 -3277 -3687 -3274
rect -3679 -3277 -3677 -3274
rect -3661 -3277 -3659 -3274
rect -3651 -3277 -3649 -3274
rect -3510 -3275 -3508 -3261
rect -3468 -3263 -3466 -3260
rect -3294 -3257 -3292 -3252
rect -3252 -3256 -3250 -3241
rect -3337 -3263 -3335 -3260
rect -3191 -3259 -3189 -3238
rect -3170 -3242 -3168 -3238
rect -3170 -3259 -3168 -3256
rect -3407 -3266 -3405 -3263
rect -3386 -3279 -3384 -3263
rect -3294 -3275 -3292 -3261
rect -3252 -3263 -3250 -3260
rect -3191 -3266 -3189 -3263
rect -3170 -3279 -3168 -3263
rect -3728 -3283 -3726 -3280
rect -4289 -3349 -4287 -3346
rect -3797 -3377 -3795 -3374
rect -3758 -3381 -3756 -3378
rect -3748 -3381 -3746 -3378
rect -5090 -3399 -5088 -3396
rect -6072 -3452 -6070 -3449
rect -6033 -3456 -6031 -3453
rect -6023 -3456 -6021 -3453
rect -6072 -3478 -6070 -3464
rect -6005 -3462 -6003 -3459
rect -5995 -3462 -5993 -3459
rect -6072 -3487 -6070 -3484
rect -6033 -3489 -6031 -3480
rect -6023 -3490 -6021 -3480
rect -6072 -3507 -6070 -3504
rect -6072 -3533 -6070 -3519
rect -6033 -3521 -6031 -3494
rect -6023 -3521 -6021 -3495
rect -6005 -3497 -6003 -3486
rect -6005 -3521 -6003 -3501
rect -5995 -3508 -5993 -3486
rect -4289 -3407 -4287 -3389
rect -3797 -3403 -3795 -3389
rect -3730 -3387 -3728 -3384
rect -3720 -3387 -3718 -3384
rect -3797 -3412 -3795 -3409
rect -3758 -3414 -3756 -3405
rect -3748 -3415 -3746 -3405
rect -4289 -3431 -4287 -3427
rect -3797 -3432 -3795 -3429
rect -3797 -3458 -3795 -3444
rect -3758 -3446 -3756 -3419
rect -3748 -3446 -3746 -3420
rect -3730 -3422 -3728 -3411
rect -3730 -3446 -3728 -3426
rect -3720 -3433 -3718 -3411
rect -3515 -3415 -3513 -3398
rect -3412 -3413 -3410 -3411
rect -3391 -3414 -3389 -3395
rect -3299 -3415 -3297 -3398
rect -3196 -3413 -3194 -3411
rect -3175 -3414 -3173 -3395
rect -3720 -3446 -3718 -3437
rect -3558 -3440 -3556 -3425
rect -3515 -3432 -3513 -3425
rect -3515 -3441 -3513 -3436
rect -3473 -3440 -3471 -3425
rect -3558 -3447 -3556 -3444
rect -3412 -3443 -3410 -3422
rect -3391 -3426 -3389 -3422
rect -3342 -3440 -3340 -3425
rect -3299 -3432 -3297 -3425
rect -3391 -3443 -3389 -3440
rect -3758 -3461 -3756 -3458
rect -3748 -3461 -3746 -3458
rect -3730 -3461 -3728 -3458
rect -3720 -3461 -3718 -3458
rect -3515 -3459 -3513 -3445
rect -3473 -3447 -3471 -3444
rect -3299 -3441 -3297 -3436
rect -3257 -3440 -3255 -3425
rect -3342 -3447 -3340 -3444
rect -3196 -3443 -3194 -3422
rect -3175 -3426 -3173 -3422
rect -3175 -3443 -3173 -3440
rect -3412 -3450 -3410 -3447
rect -3391 -3463 -3389 -3447
rect -3299 -3459 -3297 -3445
rect -3257 -3447 -3255 -3444
rect -3196 -3450 -3194 -3447
rect -3175 -3463 -3173 -3447
rect -3797 -3467 -3795 -3464
rect -4288 -3480 -4286 -3477
rect -4918 -3488 -4916 -3485
rect -5995 -3521 -5993 -3512
rect -5090 -3515 -5088 -3499
rect -6033 -3536 -6031 -3533
rect -6023 -3536 -6021 -3533
rect -6005 -3536 -6003 -3533
rect -5995 -3536 -5993 -3533
rect -6072 -3542 -6070 -3539
rect -3802 -3507 -3800 -3504
rect -3763 -3511 -3761 -3508
rect -3753 -3511 -3751 -3508
rect -4288 -3538 -4286 -3520
rect -3802 -3533 -3800 -3519
rect -3735 -3517 -3733 -3514
rect -3725 -3517 -3723 -3514
rect -3802 -3542 -3800 -3539
rect -3763 -3544 -3761 -3535
rect -3753 -3545 -3751 -3535
rect -4288 -3562 -4286 -3558
rect -3802 -3562 -3800 -3559
rect -3802 -3588 -3800 -3574
rect -3763 -3576 -3761 -3549
rect -3753 -3576 -3751 -3550
rect -3735 -3552 -3733 -3541
rect -3735 -3576 -3733 -3556
rect -3725 -3563 -3723 -3541
rect -3518 -3546 -3516 -3529
rect -3415 -3544 -3413 -3542
rect -3394 -3545 -3392 -3526
rect -3302 -3546 -3300 -3529
rect -3199 -3544 -3197 -3542
rect -3178 -3545 -3176 -3526
rect -3725 -3576 -3723 -3567
rect -3561 -3571 -3559 -3556
rect -3518 -3563 -3516 -3556
rect -3518 -3572 -3516 -3567
rect -3476 -3571 -3474 -3556
rect -3561 -3578 -3559 -3575
rect -3415 -3574 -3413 -3553
rect -3394 -3557 -3392 -3553
rect -3345 -3571 -3343 -3556
rect -3302 -3563 -3300 -3556
rect -3394 -3574 -3392 -3571
rect -4918 -3604 -4916 -3588
rect -3763 -3591 -3761 -3588
rect -3753 -3591 -3751 -3588
rect -3735 -3591 -3733 -3588
rect -3725 -3591 -3723 -3588
rect -3518 -3590 -3516 -3576
rect -3476 -3578 -3474 -3575
rect -3302 -3572 -3300 -3567
rect -3260 -3571 -3258 -3556
rect -3345 -3578 -3343 -3575
rect -3199 -3574 -3197 -3553
rect -3178 -3557 -3176 -3553
rect -3178 -3574 -3176 -3571
rect -3415 -3581 -3413 -3578
rect -3394 -3594 -3392 -3578
rect -3302 -3590 -3300 -3576
rect -3260 -3578 -3258 -3575
rect -3199 -3581 -3197 -3578
rect -3178 -3594 -3176 -3578
rect -3802 -3597 -3800 -3594
rect -4288 -3611 -4286 -3608
rect -6079 -3624 -6077 -3621
rect -6040 -3628 -6038 -3625
rect -6030 -3628 -6028 -3625
rect -6079 -3650 -6077 -3636
rect -6012 -3634 -6010 -3631
rect -6002 -3634 -6000 -3631
rect -6079 -3659 -6077 -3656
rect -6040 -3661 -6038 -3652
rect -6030 -3662 -6028 -3652
rect -3798 -3635 -3796 -3632
rect -3759 -3639 -3757 -3636
rect -3749 -3639 -3747 -3636
rect -6079 -3679 -6077 -3676
rect -6079 -3705 -6077 -3691
rect -6040 -3693 -6038 -3666
rect -6030 -3693 -6028 -3667
rect -6012 -3669 -6010 -3658
rect -6012 -3693 -6010 -3673
rect -6002 -3680 -6000 -3658
rect -5082 -3667 -5080 -3664
rect -6002 -3693 -6000 -3684
rect -6040 -3708 -6038 -3705
rect -6030 -3708 -6028 -3705
rect -6012 -3708 -6010 -3705
rect -6002 -3708 -6000 -3705
rect -6079 -3714 -6077 -3711
rect -6076 -3768 -6074 -3765
rect -4288 -3669 -4286 -3651
rect -3798 -3661 -3796 -3647
rect -3731 -3645 -3729 -3642
rect -3721 -3645 -3719 -3642
rect -3798 -3670 -3796 -3667
rect -3759 -3672 -3757 -3663
rect -3749 -3673 -3747 -3663
rect -4288 -3693 -4286 -3689
rect -3798 -3690 -3796 -3687
rect -3798 -3716 -3796 -3702
rect -3759 -3704 -3757 -3677
rect -3749 -3704 -3747 -3678
rect -3731 -3680 -3729 -3669
rect -3731 -3704 -3729 -3684
rect -3721 -3691 -3719 -3669
rect -3531 -3676 -3529 -3659
rect -3428 -3674 -3426 -3672
rect -3407 -3675 -3405 -3656
rect -3315 -3676 -3313 -3659
rect -3212 -3674 -3210 -3672
rect -3191 -3675 -3189 -3656
rect -3721 -3704 -3719 -3695
rect -3574 -3701 -3572 -3686
rect -3531 -3693 -3529 -3686
rect -3531 -3702 -3529 -3697
rect -3489 -3701 -3487 -3686
rect -3574 -3708 -3572 -3705
rect -3428 -3704 -3426 -3683
rect -3407 -3687 -3405 -3683
rect -3358 -3701 -3356 -3686
rect -3315 -3693 -3313 -3686
rect -3407 -3704 -3405 -3701
rect -4744 -3722 -4742 -3719
rect -3759 -3719 -3757 -3716
rect -3749 -3719 -3747 -3716
rect -3731 -3719 -3729 -3716
rect -3721 -3719 -3719 -3716
rect -3531 -3720 -3529 -3706
rect -3489 -3708 -3487 -3705
rect -3315 -3702 -3313 -3697
rect -3273 -3701 -3271 -3686
rect -3358 -3708 -3356 -3705
rect -3212 -3704 -3210 -3683
rect -3191 -3687 -3189 -3683
rect -3191 -3704 -3189 -3701
rect -3428 -3711 -3426 -3708
rect -6037 -3772 -6035 -3769
rect -6027 -3772 -6025 -3769
rect -6076 -3794 -6074 -3780
rect -6009 -3778 -6007 -3775
rect -5999 -3778 -5997 -3775
rect -6076 -3803 -6074 -3800
rect -6037 -3805 -6035 -3796
rect -6027 -3806 -6025 -3796
rect -5082 -3783 -5080 -3767
rect -6076 -3823 -6074 -3820
rect -6076 -3849 -6074 -3835
rect -6037 -3837 -6035 -3810
rect -6027 -3837 -6025 -3811
rect -6009 -3813 -6007 -3802
rect -6009 -3837 -6007 -3817
rect -5999 -3824 -5997 -3802
rect -3798 -3725 -3796 -3722
rect -3407 -3724 -3405 -3708
rect -3315 -3720 -3313 -3706
rect -3273 -3708 -3271 -3705
rect -3212 -3711 -3210 -3708
rect -3191 -3724 -3189 -3708
rect -4620 -3753 -4618 -3750
rect -5999 -3837 -5997 -3828
rect -4744 -3838 -4742 -3822
rect -6037 -3852 -6035 -3849
rect -6027 -3852 -6025 -3849
rect -6009 -3852 -6007 -3849
rect -5999 -3852 -5997 -3849
rect -4289 -3754 -4287 -3751
rect -3797 -3778 -3795 -3775
rect -3758 -3782 -3756 -3779
rect -3748 -3782 -3746 -3779
rect -4289 -3812 -4287 -3794
rect -3797 -3804 -3795 -3790
rect -3730 -3788 -3728 -3785
rect -3720 -3788 -3718 -3785
rect -3797 -3813 -3795 -3810
rect -3758 -3815 -3756 -3806
rect -3748 -3816 -3746 -3806
rect -4289 -3836 -4287 -3832
rect -3797 -3833 -3795 -3830
rect -6076 -3858 -6074 -3855
rect -4620 -3869 -4618 -3853
rect -3797 -3859 -3795 -3845
rect -3758 -3847 -3756 -3820
rect -3748 -3847 -3746 -3821
rect -3730 -3823 -3728 -3812
rect -3730 -3847 -3728 -3827
rect -3720 -3834 -3718 -3812
rect -3530 -3819 -3528 -3802
rect -3427 -3817 -3425 -3815
rect -3406 -3818 -3404 -3799
rect -3314 -3819 -3312 -3802
rect -3211 -3817 -3209 -3815
rect -3190 -3818 -3188 -3799
rect -3720 -3847 -3718 -3838
rect -3573 -3844 -3571 -3829
rect -3530 -3836 -3528 -3829
rect -3530 -3845 -3528 -3840
rect -3488 -3844 -3486 -3829
rect -3573 -3851 -3571 -3848
rect -3427 -3847 -3425 -3826
rect -3406 -3830 -3404 -3826
rect -3357 -3844 -3355 -3829
rect -3314 -3836 -3312 -3829
rect -3406 -3847 -3404 -3844
rect -3758 -3862 -3756 -3859
rect -3748 -3862 -3746 -3859
rect -3730 -3862 -3728 -3859
rect -3720 -3862 -3718 -3859
rect -3530 -3863 -3528 -3849
rect -3488 -3851 -3486 -3848
rect -3314 -3845 -3312 -3840
rect -3272 -3844 -3270 -3829
rect -3357 -3851 -3355 -3848
rect -3211 -3847 -3209 -3826
rect -3190 -3830 -3188 -3826
rect -3190 -3847 -3188 -3844
rect -3427 -3854 -3425 -3851
rect -3797 -3868 -3795 -3865
rect -3406 -3867 -3404 -3851
rect -3314 -3863 -3312 -3849
rect -3272 -3851 -3270 -3848
rect -3211 -3854 -3209 -3851
rect -3190 -3867 -3188 -3851
rect -4289 -3906 -4287 -3903
rect -6080 -3916 -6078 -3913
rect -4480 -3916 -4478 -3913
rect -6041 -3920 -6039 -3917
rect -6031 -3920 -6029 -3917
rect -6080 -3942 -6078 -3928
rect -6013 -3926 -6011 -3923
rect -6003 -3926 -6001 -3923
rect -6080 -3951 -6078 -3948
rect -6041 -3953 -6039 -3944
rect -6031 -3954 -6029 -3944
rect -6080 -3971 -6078 -3968
rect -6080 -3997 -6078 -3983
rect -6041 -3985 -6039 -3958
rect -6031 -3985 -6029 -3959
rect -6013 -3961 -6011 -3950
rect -6013 -3985 -6011 -3965
rect -6003 -3972 -6001 -3950
rect -6003 -3985 -6001 -3976
rect -6041 -4000 -6039 -3997
rect -6031 -4000 -6029 -3997
rect -6013 -4000 -6011 -3997
rect -6003 -4000 -6001 -3997
rect -6080 -4006 -6078 -4003
rect -3545 -3937 -3543 -3920
rect -3442 -3935 -3440 -3933
rect -3421 -3936 -3419 -3917
rect -4289 -3964 -4287 -3946
rect -3329 -3937 -3327 -3920
rect -3226 -3935 -3224 -3933
rect -3205 -3936 -3203 -3917
rect -3588 -3962 -3586 -3947
rect -3545 -3954 -3543 -3947
rect -3545 -3963 -3543 -3958
rect -3503 -3962 -3501 -3947
rect -3588 -3969 -3586 -3966
rect -3442 -3965 -3440 -3944
rect -3421 -3948 -3419 -3944
rect -3372 -3962 -3370 -3947
rect -3329 -3954 -3327 -3947
rect -3421 -3965 -3419 -3962
rect -3545 -3981 -3543 -3967
rect -3503 -3969 -3501 -3966
rect -3329 -3963 -3327 -3958
rect -3287 -3962 -3285 -3947
rect -3372 -3969 -3370 -3966
rect -3226 -3965 -3224 -3944
rect -3205 -3948 -3203 -3944
rect -3205 -3965 -3203 -3962
rect -3442 -3972 -3440 -3969
rect -4289 -3988 -4287 -3984
rect -3421 -3985 -3419 -3969
rect -3329 -3981 -3327 -3967
rect -3287 -3969 -3285 -3966
rect -3226 -3972 -3224 -3969
rect -3205 -3985 -3203 -3969
rect -4480 -4032 -4478 -4016
rect -6055 -4132 -6053 -4129
rect -6016 -4136 -6014 -4133
rect -6006 -4136 -6004 -4133
rect -6055 -4158 -6053 -4144
rect -5988 -4142 -5986 -4139
rect -5978 -4142 -5976 -4139
rect -6055 -4167 -6053 -4164
rect -6016 -4169 -6014 -4160
rect -6006 -4170 -6004 -4160
rect -6055 -4187 -6053 -4184
rect -6055 -4213 -6053 -4199
rect -6016 -4201 -6014 -4174
rect -6006 -4201 -6004 -4175
rect -5988 -4177 -5986 -4166
rect -5988 -4201 -5986 -4181
rect -5978 -4188 -5976 -4166
rect -5978 -4201 -5976 -4192
rect -6016 -4216 -6014 -4213
rect -6006 -4216 -6004 -4213
rect -5988 -4216 -5986 -4213
rect -5978 -4216 -5976 -4213
rect -6055 -4222 -6053 -4219
rect -4909 -4291 -4907 -4288
rect -6056 -4375 -6054 -4372
rect -6045 -4375 -6043 -4372
rect -6014 -4382 -6012 -4378
rect -6056 -4424 -6054 -4395
rect -6045 -4424 -6043 -4395
rect -4735 -4324 -4733 -4321
rect -6014 -4416 -6012 -4402
rect -4909 -4407 -4907 -4391
rect -4611 -4395 -4609 -4392
rect -6014 -4429 -6012 -4426
rect -4735 -4440 -4733 -4424
rect -6056 -4447 -6054 -4444
rect -6045 -4447 -6043 -4444
rect -6055 -4484 -6053 -4481
rect -6044 -4484 -6042 -4481
rect -6013 -4491 -6011 -4487
rect -6055 -4533 -6053 -4504
rect -6044 -4533 -6042 -4504
rect -4472 -4494 -4470 -4491
rect -4611 -4511 -4609 -4495
rect -6013 -4525 -6011 -4511
rect -6013 -4538 -6011 -4535
rect -6055 -4556 -6053 -4553
rect -6044 -4556 -6042 -4553
rect -4393 -4553 -4391 -4550
rect -6052 -4612 -6050 -4609
rect -6041 -4612 -6039 -4609
rect -4472 -4610 -4470 -4594
rect -6010 -4619 -6008 -4615
rect -6052 -4661 -6050 -4632
rect -6041 -4661 -6039 -4632
rect -6010 -4653 -6008 -4639
rect -6010 -4666 -6008 -4663
rect -4393 -4669 -4391 -4653
rect -6052 -4684 -6050 -4681
rect -6041 -4684 -6039 -4681
rect -6050 -4732 -6048 -4729
rect -6039 -4732 -6037 -4729
rect -6008 -4739 -6006 -4735
rect -6050 -4781 -6048 -4752
rect -6039 -4781 -6037 -4752
rect -6008 -4773 -6006 -4759
rect -6008 -4786 -6006 -4783
rect -6050 -4804 -6048 -4801
rect -6039 -4804 -6037 -4801
rect -5073 -4811 -5071 -4808
rect -6048 -4873 -6046 -4870
rect -6037 -4873 -6035 -4870
rect -5226 -4872 -5224 -4869
rect -6006 -4880 -6004 -4876
rect -6048 -4922 -6046 -4893
rect -6037 -4922 -6035 -4893
rect -6006 -4914 -6004 -4900
rect -6006 -4927 -6004 -4924
rect -5226 -4930 -5224 -4912
rect -5073 -4927 -5071 -4911
rect -6048 -4945 -6046 -4942
rect -6037 -4945 -6035 -4942
rect -5226 -4954 -5224 -4950
<< polycontact >>
rect -7704 -2628 -7700 -2624
rect -8122 -2634 -8118 -2630
rect -7980 -2637 -7976 -2633
rect -7838 -2635 -7834 -2631
rect -7569 -2634 -7565 -2630
rect -7449 -2633 -7445 -2629
rect -7329 -2633 -7325 -2629
rect -7204 -2632 -7200 -2628
rect -7086 -2632 -7082 -2628
rect -6967 -2630 -6963 -2626
rect -7726 -2671 -7722 -2667
rect -7669 -2671 -7665 -2667
rect -8144 -2677 -8140 -2673
rect -8087 -2677 -8083 -2673
rect -8002 -2680 -7998 -2676
rect -7945 -2680 -7941 -2676
rect -7860 -2678 -7856 -2674
rect -7803 -2678 -7799 -2674
rect -7591 -2677 -7587 -2673
rect -7534 -2677 -7530 -2673
rect -7471 -2676 -7467 -2672
rect -7414 -2676 -7410 -2672
rect -7351 -2676 -7347 -2672
rect -7294 -2676 -7290 -2672
rect -7226 -2675 -7222 -2671
rect -7169 -2675 -7165 -2671
rect -7108 -2675 -7104 -2671
rect -7051 -2675 -7047 -2671
rect -6989 -2673 -6985 -2669
rect -6932 -2673 -6928 -2669
rect -7704 -2713 -7700 -2709
rect -8122 -2719 -8118 -2715
rect -7980 -2722 -7976 -2718
rect -7838 -2720 -7834 -2716
rect -7569 -2719 -7565 -2715
rect -7449 -2718 -7445 -2714
rect -7329 -2718 -7325 -2714
rect -7204 -2717 -7200 -2713
rect -7086 -2717 -7082 -2713
rect -6967 -2715 -6963 -2711
rect -7704 -2774 -7700 -2770
rect -8122 -2780 -8118 -2776
rect -7980 -2783 -7976 -2779
rect -7838 -2781 -7834 -2777
rect -7569 -2780 -7565 -2776
rect -7449 -2779 -7445 -2775
rect -7329 -2779 -7325 -2775
rect -7204 -2778 -7200 -2774
rect -7086 -2778 -7082 -2774
rect -6967 -2776 -6963 -2772
rect -7730 -2795 -7726 -2791
rect -7666 -2795 -7662 -2791
rect -8148 -2801 -8144 -2797
rect -8084 -2801 -8080 -2797
rect -8006 -2804 -8002 -2800
rect -7942 -2804 -7938 -2800
rect -7864 -2802 -7860 -2798
rect -7800 -2802 -7796 -2798
rect -7595 -2801 -7591 -2797
rect -7531 -2801 -7527 -2797
rect -7475 -2800 -7471 -2796
rect -7411 -2800 -7407 -2796
rect -7355 -2800 -7351 -2796
rect -7291 -2800 -7287 -2796
rect -7230 -2799 -7226 -2795
rect -7166 -2799 -7162 -2795
rect -7112 -2799 -7108 -2795
rect -7048 -2799 -7044 -2795
rect -6993 -2797 -6989 -2793
rect -6929 -2797 -6925 -2793
rect -7704 -2844 -7700 -2840
rect -8122 -2850 -8118 -2846
rect -7980 -2853 -7976 -2849
rect -7838 -2851 -7834 -2847
rect -7569 -2850 -7565 -2846
rect -7449 -2849 -7445 -2845
rect -7329 -2849 -7325 -2845
rect -7204 -2848 -7200 -2844
rect -7086 -2848 -7082 -2844
rect -6967 -2846 -6963 -2842
rect -7726 -2887 -7722 -2883
rect -7669 -2887 -7665 -2883
rect -8144 -2893 -8140 -2889
rect -8087 -2893 -8083 -2889
rect -8002 -2896 -7998 -2892
rect -7945 -2896 -7941 -2892
rect -7860 -2894 -7856 -2890
rect -7803 -2894 -7799 -2890
rect -7591 -2893 -7587 -2889
rect -7534 -2893 -7530 -2889
rect -7471 -2892 -7467 -2888
rect -7414 -2892 -7410 -2888
rect -7351 -2892 -7347 -2888
rect -7294 -2892 -7290 -2888
rect -7226 -2891 -7222 -2887
rect -7169 -2891 -7165 -2887
rect -7108 -2891 -7104 -2887
rect -7051 -2891 -7047 -2887
rect -6989 -2889 -6985 -2885
rect -6932 -2889 -6928 -2885
rect -7704 -2929 -7700 -2925
rect -8122 -2935 -8118 -2931
rect -7980 -2938 -7976 -2934
rect -7838 -2936 -7834 -2932
rect -7569 -2935 -7565 -2931
rect -7449 -2934 -7445 -2930
rect -7329 -2934 -7325 -2930
rect -7204 -2933 -7200 -2929
rect -7086 -2933 -7082 -2929
rect -6967 -2931 -6963 -2927
rect -7704 -2990 -7700 -2986
rect -8122 -2996 -8118 -2992
rect -7980 -2999 -7976 -2995
rect -7838 -2997 -7834 -2993
rect -7569 -2996 -7565 -2992
rect -7449 -2995 -7445 -2991
rect -7329 -2995 -7325 -2991
rect -7204 -2994 -7200 -2990
rect -7086 -2994 -7082 -2990
rect -6967 -2992 -6963 -2988
rect -7730 -3011 -7726 -3007
rect -7666 -3011 -7662 -3007
rect -8148 -3017 -8144 -3013
rect -8084 -3017 -8080 -3013
rect -8006 -3020 -8002 -3016
rect -7942 -3020 -7938 -3016
rect -7864 -3018 -7860 -3014
rect -7800 -3018 -7796 -3014
rect -7595 -3017 -7591 -3013
rect -7531 -3017 -7527 -3013
rect -7475 -3016 -7471 -3012
rect -7411 -3016 -7407 -3012
rect -7355 -3016 -7351 -3012
rect -7291 -3016 -7287 -3012
rect -7230 -3015 -7226 -3011
rect -7166 -3015 -7162 -3011
rect -7112 -3015 -7108 -3011
rect -7048 -3015 -7044 -3011
rect -6993 -3013 -6989 -3009
rect -6929 -3013 -6925 -3009
rect -3732 -3216 -3728 -3212
rect -3514 -3218 -3510 -3214
rect -3732 -3271 -3728 -3267
rect -3663 -3242 -3659 -3238
rect -3390 -3215 -3386 -3211
rect -3298 -3218 -3294 -3214
rect -3174 -3215 -3170 -3211
rect -3652 -3253 -3648 -3249
rect -3557 -3253 -3553 -3249
rect -3472 -3253 -3468 -3249
rect -3411 -3253 -3407 -3249
rect -3341 -3253 -3337 -3249
rect -3514 -3275 -3510 -3271
rect -3256 -3253 -3252 -3249
rect -3195 -3253 -3191 -3249
rect -3390 -3279 -3386 -3275
rect -3298 -3275 -3294 -3271
rect -3174 -3279 -3170 -3275
rect -6076 -3475 -6072 -3471
rect -6076 -3530 -6072 -3526
rect -6007 -3501 -6003 -3497
rect -3801 -3400 -3797 -3396
rect -3519 -3402 -3515 -3398
rect -3801 -3455 -3797 -3451
rect -3732 -3426 -3728 -3422
rect -3395 -3399 -3391 -3395
rect -3303 -3402 -3299 -3398
rect -3179 -3399 -3175 -3395
rect -3721 -3437 -3717 -3433
rect -3562 -3437 -3558 -3433
rect -3477 -3437 -3473 -3433
rect -3416 -3437 -3412 -3433
rect -3346 -3437 -3342 -3433
rect -3519 -3459 -3515 -3455
rect -3261 -3437 -3257 -3433
rect -3200 -3437 -3196 -3433
rect -3395 -3463 -3391 -3459
rect -3303 -3459 -3299 -3455
rect -3179 -3463 -3175 -3459
rect -5996 -3512 -5992 -3508
rect -3806 -3530 -3802 -3526
rect -3522 -3533 -3518 -3529
rect -3806 -3585 -3802 -3581
rect -3737 -3556 -3733 -3552
rect -3398 -3530 -3394 -3526
rect -3306 -3533 -3302 -3529
rect -3182 -3530 -3178 -3526
rect -3726 -3567 -3722 -3563
rect -3565 -3568 -3561 -3564
rect -3480 -3568 -3476 -3564
rect -3419 -3568 -3415 -3564
rect -3349 -3568 -3345 -3564
rect -3522 -3590 -3518 -3586
rect -3264 -3568 -3260 -3564
rect -3203 -3568 -3199 -3564
rect -3398 -3594 -3394 -3590
rect -3306 -3590 -3302 -3586
rect -3182 -3594 -3178 -3590
rect -6083 -3647 -6079 -3643
rect -6083 -3702 -6079 -3698
rect -6014 -3673 -6010 -3669
rect -6003 -3684 -5999 -3680
rect -3802 -3658 -3798 -3654
rect -3535 -3663 -3531 -3659
rect -3802 -3713 -3798 -3709
rect -3733 -3684 -3729 -3680
rect -3411 -3660 -3407 -3656
rect -3319 -3663 -3315 -3659
rect -3195 -3660 -3191 -3656
rect -3722 -3695 -3718 -3691
rect -3578 -3698 -3574 -3694
rect -3493 -3698 -3489 -3694
rect -3432 -3698 -3428 -3694
rect -3362 -3698 -3358 -3694
rect -3535 -3720 -3531 -3716
rect -3277 -3698 -3273 -3694
rect -3216 -3698 -3212 -3694
rect -6080 -3791 -6076 -3787
rect -6080 -3846 -6076 -3842
rect -6011 -3817 -6007 -3813
rect -3411 -3724 -3407 -3720
rect -3319 -3720 -3315 -3716
rect -3195 -3724 -3191 -3720
rect -6000 -3828 -5996 -3824
rect -3801 -3801 -3797 -3797
rect -3534 -3806 -3530 -3802
rect -3801 -3856 -3797 -3852
rect -3732 -3827 -3728 -3823
rect -3410 -3803 -3406 -3799
rect -3318 -3806 -3314 -3802
rect -3194 -3803 -3190 -3799
rect -3721 -3838 -3717 -3834
rect -3577 -3841 -3573 -3837
rect -3492 -3841 -3488 -3837
rect -3431 -3841 -3427 -3837
rect -3361 -3841 -3357 -3837
rect -3534 -3863 -3530 -3859
rect -3276 -3841 -3272 -3837
rect -3215 -3841 -3211 -3837
rect -3410 -3867 -3406 -3863
rect -3318 -3863 -3314 -3859
rect -3194 -3867 -3190 -3863
rect -6084 -3939 -6080 -3935
rect -6084 -3994 -6080 -3990
rect -6015 -3965 -6011 -3961
rect -6004 -3976 -6000 -3972
rect -3549 -3924 -3545 -3920
rect -3425 -3921 -3421 -3917
rect -3333 -3924 -3329 -3920
rect -3209 -3921 -3205 -3917
rect -3592 -3959 -3588 -3955
rect -3507 -3959 -3503 -3955
rect -3446 -3959 -3442 -3955
rect -3376 -3959 -3372 -3955
rect -3549 -3981 -3545 -3977
rect -3291 -3959 -3287 -3955
rect -3230 -3959 -3226 -3955
rect -3425 -3985 -3421 -3981
rect -3333 -3981 -3329 -3977
rect -3209 -3985 -3205 -3981
rect -6059 -4155 -6055 -4151
rect -6059 -4210 -6055 -4206
rect -5990 -4181 -5986 -4177
rect -5979 -4192 -5975 -4188
rect -6060 -4421 -6056 -4417
rect -6049 -4414 -6045 -4410
rect -6018 -4413 -6014 -4409
rect -6059 -4530 -6055 -4526
rect -6048 -4523 -6044 -4519
rect -6017 -4522 -6013 -4518
rect -6056 -4658 -6052 -4654
rect -6045 -4651 -6041 -4647
rect -6014 -4650 -6010 -4646
rect -6054 -4778 -6050 -4774
rect -6043 -4771 -6039 -4767
rect -6012 -4770 -6008 -4766
rect -6052 -4919 -6048 -4915
rect -6041 -4912 -6037 -4908
rect -6010 -4911 -6006 -4907
<< polypplus >>
rect -7684 -2630 -7681 -2628
rect -8102 -2636 -8099 -2634
rect -6947 -2632 -6944 -2630
rect -7818 -2637 -7815 -2635
rect -7549 -2636 -7546 -2634
rect -7429 -2635 -7426 -2633
rect -7309 -2635 -7306 -2633
rect -7184 -2634 -7181 -2632
rect -7066 -2634 -7063 -2632
rect -7960 -2639 -7957 -2637
rect -7684 -2673 -7682 -2671
rect -8102 -2679 -8100 -2677
rect -7818 -2680 -7816 -2678
rect -7549 -2679 -7547 -2677
rect -7429 -2678 -7427 -2676
rect -7309 -2678 -7307 -2676
rect -7184 -2677 -7182 -2675
rect -6947 -2675 -6945 -2673
rect -7066 -2677 -7064 -2675
rect -7960 -2682 -7958 -2680
rect -7684 -2715 -7681 -2713
rect -8102 -2721 -8099 -2719
rect -6947 -2717 -6944 -2715
rect -7818 -2722 -7815 -2720
rect -7549 -2721 -7546 -2719
rect -7429 -2720 -7426 -2718
rect -7309 -2720 -7306 -2718
rect -7184 -2719 -7181 -2717
rect -7066 -2719 -7063 -2717
rect -7960 -2724 -7957 -2722
rect -7681 -2776 -7680 -2774
rect -8099 -2782 -8098 -2780
rect -6944 -2778 -6943 -2776
rect -7815 -2783 -7814 -2781
rect -7546 -2782 -7545 -2780
rect -7426 -2781 -7425 -2779
rect -7306 -2781 -7305 -2779
rect -7181 -2780 -7180 -2778
rect -7063 -2780 -7062 -2778
rect -7957 -2785 -7956 -2783
rect -7684 -2846 -7681 -2844
rect -8102 -2852 -8099 -2850
rect -6947 -2848 -6944 -2846
rect -7818 -2853 -7815 -2851
rect -7549 -2852 -7546 -2850
rect -7429 -2851 -7426 -2849
rect -7309 -2851 -7306 -2849
rect -7184 -2850 -7181 -2848
rect -7066 -2850 -7063 -2848
rect -7960 -2855 -7957 -2853
rect -7684 -2889 -7682 -2887
rect -8102 -2895 -8100 -2893
rect -7818 -2896 -7816 -2894
rect -7549 -2895 -7547 -2893
rect -7429 -2894 -7427 -2892
rect -7309 -2894 -7307 -2892
rect -7184 -2893 -7182 -2891
rect -6947 -2891 -6945 -2889
rect -7066 -2893 -7064 -2891
rect -7960 -2898 -7958 -2896
rect -7684 -2931 -7681 -2929
rect -8102 -2937 -8099 -2935
rect -6947 -2933 -6944 -2931
rect -7818 -2938 -7815 -2936
rect -7549 -2937 -7546 -2935
rect -7429 -2936 -7426 -2934
rect -7309 -2936 -7306 -2934
rect -7184 -2935 -7181 -2933
rect -7066 -2935 -7063 -2933
rect -7960 -2940 -7957 -2938
rect -7681 -2992 -7680 -2990
rect -8099 -2998 -8098 -2996
rect -6944 -2994 -6943 -2992
rect -7815 -2999 -7814 -2997
rect -7546 -2998 -7545 -2996
rect -7426 -2997 -7425 -2995
rect -7306 -2997 -7305 -2995
rect -7181 -2996 -7180 -2994
rect -7063 -2996 -7062 -2994
rect -7957 -3001 -7956 -2999
rect -3553 -3233 -3551 -3230
rect -3407 -3230 -3405 -3229
rect -3510 -3233 -3508 -3231
rect -3468 -3233 -3466 -3230
rect -3337 -3233 -3335 -3230
rect -3191 -3230 -3189 -3229
rect -3294 -3233 -3292 -3231
rect -3252 -3233 -3250 -3230
rect -3558 -3417 -3556 -3414
rect -3412 -3414 -3410 -3413
rect -3515 -3417 -3513 -3415
rect -3473 -3417 -3471 -3414
rect -3342 -3417 -3340 -3414
rect -3196 -3414 -3194 -3413
rect -3299 -3417 -3297 -3415
rect -3257 -3417 -3255 -3414
rect -3561 -3548 -3559 -3545
rect -3415 -3545 -3413 -3544
rect -3518 -3548 -3516 -3546
rect -3476 -3548 -3474 -3545
rect -3345 -3548 -3343 -3545
rect -3199 -3545 -3197 -3544
rect -3302 -3548 -3300 -3546
rect -3260 -3548 -3258 -3545
rect -3574 -3678 -3572 -3675
rect -3428 -3675 -3426 -3674
rect -3531 -3678 -3529 -3676
rect -3489 -3678 -3487 -3675
rect -3358 -3678 -3356 -3675
rect -3212 -3675 -3210 -3674
rect -3315 -3678 -3313 -3676
rect -3273 -3678 -3271 -3675
rect -3573 -3821 -3571 -3818
rect -3427 -3818 -3425 -3817
rect -3530 -3821 -3528 -3819
rect -3488 -3821 -3486 -3818
rect -3357 -3821 -3355 -3818
rect -3211 -3818 -3209 -3817
rect -3314 -3821 -3312 -3819
rect -3272 -3821 -3270 -3818
rect -3588 -3939 -3586 -3936
rect -3442 -3936 -3440 -3935
rect -3545 -3939 -3543 -3937
rect -3503 -3939 -3501 -3936
rect -3372 -3939 -3370 -3936
rect -3226 -3936 -3224 -3935
rect -3329 -3939 -3327 -3937
rect -3287 -3939 -3285 -3936
<< metal1 >>
rect -8136 -2629 -8133 -2623
rect -8136 -2633 -8129 -2629
rect -8122 -2630 -8118 -2612
rect -8098 -2629 -8094 -2623
rect -8136 -2648 -8133 -2633
rect -8102 -2633 -8094 -2629
rect -8125 -2641 -8110 -2637
rect -8147 -2663 -8140 -2659
rect -8144 -2673 -8140 -2663
rect -8122 -2672 -8118 -2641
rect -8098 -2648 -8094 -2633
rect -7994 -2632 -7991 -2626
rect -7994 -2636 -7987 -2632
rect -7980 -2633 -7976 -2615
rect -7956 -2632 -7952 -2626
rect -7994 -2651 -7991 -2636
rect -7960 -2636 -7952 -2632
rect -7983 -2644 -7968 -2640
rect -8126 -2676 -8110 -2672
rect -8087 -2673 -8083 -2661
rect -8005 -2666 -7998 -2662
rect -8002 -2676 -7998 -2666
rect -7980 -2675 -7976 -2644
rect -7956 -2651 -7952 -2636
rect -7852 -2630 -7849 -2624
rect -7852 -2634 -7845 -2630
rect -7838 -2631 -7834 -2613
rect -7718 -2623 -7715 -2617
rect -7814 -2630 -7810 -2624
rect -7852 -2649 -7849 -2634
rect -7818 -2634 -7810 -2630
rect -7841 -2642 -7826 -2638
rect -7863 -2664 -7856 -2660
rect -7984 -2679 -7968 -2675
rect -7945 -2676 -7941 -2664
rect -7860 -2674 -7856 -2664
rect -7838 -2673 -7834 -2642
rect -7814 -2649 -7810 -2634
rect -7718 -2627 -7711 -2623
rect -7704 -2624 -7700 -2606
rect -7680 -2623 -7676 -2617
rect -7718 -2642 -7715 -2627
rect -7684 -2627 -7676 -2623
rect -7707 -2635 -7692 -2631
rect -7729 -2657 -7722 -2653
rect -7842 -2677 -7826 -2673
rect -7803 -2674 -7799 -2662
rect -7726 -2667 -7722 -2657
rect -7704 -2666 -7700 -2635
rect -7680 -2642 -7676 -2627
rect -7583 -2629 -7580 -2623
rect -7583 -2633 -7576 -2629
rect -7569 -2630 -7565 -2612
rect -7545 -2629 -7541 -2623
rect -7583 -2648 -7580 -2633
rect -7549 -2633 -7541 -2629
rect -7572 -2641 -7557 -2637
rect -7708 -2670 -7692 -2666
rect -7669 -2667 -7665 -2655
rect -7594 -2663 -7587 -2659
rect -7591 -2673 -7587 -2663
rect -7569 -2672 -7565 -2641
rect -7545 -2648 -7541 -2633
rect -7463 -2628 -7460 -2622
rect -7463 -2632 -7456 -2628
rect -7449 -2629 -7445 -2611
rect -7425 -2628 -7421 -2622
rect -7463 -2647 -7460 -2632
rect -7429 -2632 -7421 -2628
rect -7452 -2640 -7437 -2636
rect -7708 -2678 -7692 -2674
rect -7573 -2676 -7557 -2672
rect -7534 -2673 -7530 -2661
rect -7474 -2662 -7467 -2658
rect -7471 -2672 -7467 -2662
rect -7449 -2671 -7445 -2640
rect -7425 -2647 -7421 -2632
rect -7343 -2628 -7340 -2622
rect -7343 -2632 -7336 -2628
rect -7329 -2629 -7325 -2611
rect -7305 -2628 -7301 -2622
rect -7343 -2647 -7340 -2632
rect -7309 -2632 -7301 -2628
rect -7332 -2640 -7317 -2636
rect -7453 -2675 -7437 -2671
rect -7414 -2672 -7410 -2660
rect -7354 -2662 -7347 -2658
rect -7351 -2672 -7347 -2662
rect -7329 -2671 -7325 -2640
rect -7305 -2647 -7301 -2632
rect -7218 -2627 -7215 -2621
rect -7218 -2631 -7211 -2627
rect -7204 -2628 -7200 -2610
rect -7180 -2627 -7176 -2621
rect -7218 -2646 -7215 -2631
rect -7184 -2631 -7176 -2627
rect -7207 -2639 -7192 -2635
rect -7333 -2675 -7317 -2671
rect -7294 -2672 -7290 -2660
rect -7229 -2661 -7222 -2657
rect -7226 -2671 -7222 -2661
rect -7204 -2670 -7200 -2639
rect -7180 -2646 -7176 -2631
rect -7100 -2627 -7097 -2621
rect -7100 -2631 -7093 -2627
rect -7086 -2628 -7082 -2610
rect -7062 -2627 -7058 -2621
rect -7100 -2646 -7097 -2631
rect -7066 -2631 -7058 -2627
rect -7089 -2639 -7074 -2635
rect -7208 -2674 -7192 -2670
rect -7169 -2671 -7165 -2659
rect -7111 -2661 -7104 -2657
rect -7108 -2671 -7104 -2661
rect -7086 -2670 -7082 -2639
rect -7062 -2646 -7058 -2631
rect -6981 -2625 -6978 -2619
rect -6981 -2629 -6974 -2625
rect -6967 -2626 -6963 -2608
rect -6943 -2625 -6939 -2619
rect -6981 -2644 -6978 -2629
rect -6947 -2629 -6939 -2625
rect -6970 -2637 -6955 -2633
rect -6992 -2659 -6985 -2655
rect -7090 -2674 -7074 -2670
rect -7051 -2671 -7047 -2659
rect -6989 -2669 -6985 -2659
rect -6967 -2668 -6963 -2637
rect -6943 -2644 -6939 -2629
rect -6971 -2672 -6955 -2668
rect -6932 -2669 -6928 -2657
rect -8126 -2684 -8110 -2680
rect -8136 -2714 -8133 -2708
rect -8136 -2718 -8129 -2714
rect -8122 -2715 -8118 -2684
rect -7984 -2687 -7968 -2683
rect -7842 -2685 -7826 -2681
rect -8098 -2714 -8094 -2708
rect -8136 -2733 -8133 -2718
rect -8102 -2718 -8094 -2714
rect -8125 -2726 -8110 -2722
rect -8141 -2779 -8132 -2775
rect -8122 -2776 -8118 -2726
rect -8098 -2733 -8094 -2718
rect -7994 -2717 -7991 -2711
rect -7994 -2721 -7987 -2717
rect -7980 -2718 -7976 -2687
rect -7956 -2717 -7952 -2711
rect -7994 -2736 -7991 -2721
rect -7960 -2721 -7952 -2717
rect -7983 -2729 -7968 -2725
rect -8148 -2797 -8144 -2788
rect -8141 -2796 -8137 -2779
rect -8099 -2779 -8091 -2775
rect -8128 -2787 -8107 -2783
rect -8141 -2800 -8132 -2796
rect -8141 -2808 -8132 -2804
rect -8141 -2817 -8137 -2808
rect -8136 -2845 -8133 -2839
rect -8136 -2849 -8129 -2845
rect -8122 -2846 -8118 -2787
rect -8095 -2796 -8091 -2779
rect -7999 -2782 -7990 -2778
rect -7980 -2779 -7976 -2729
rect -7956 -2736 -7952 -2721
rect -7852 -2715 -7849 -2709
rect -7852 -2719 -7845 -2715
rect -7838 -2716 -7834 -2685
rect -7718 -2708 -7715 -2702
rect -7814 -2715 -7810 -2709
rect -7852 -2734 -7849 -2719
rect -7818 -2719 -7810 -2715
rect -7841 -2727 -7826 -2723
rect -8099 -2800 -8091 -2796
rect -8084 -2797 -8080 -2787
rect -8006 -2800 -8002 -2791
rect -7999 -2799 -7995 -2782
rect -7957 -2782 -7949 -2778
rect -7986 -2790 -7965 -2786
rect -7999 -2803 -7990 -2799
rect -8099 -2808 -8091 -2804
rect -8095 -2817 -8091 -2808
rect -7999 -2811 -7990 -2807
rect -7999 -2820 -7995 -2811
rect -8098 -2845 -8094 -2839
rect -8136 -2864 -8133 -2849
rect -8102 -2849 -8094 -2845
rect -8125 -2857 -8110 -2853
rect -8144 -2889 -8140 -2875
rect -8122 -2888 -8118 -2857
rect -8098 -2864 -8094 -2849
rect -7994 -2848 -7991 -2842
rect -7994 -2852 -7987 -2848
rect -7980 -2849 -7976 -2790
rect -7953 -2799 -7949 -2782
rect -7857 -2780 -7848 -2776
rect -7838 -2777 -7834 -2727
rect -7814 -2734 -7810 -2719
rect -7718 -2712 -7711 -2708
rect -7704 -2709 -7700 -2678
rect -7573 -2684 -7557 -2680
rect -7453 -2683 -7437 -2679
rect -7333 -2683 -7317 -2679
rect -7208 -2682 -7192 -2678
rect -7090 -2682 -7074 -2678
rect -6971 -2680 -6955 -2676
rect -7680 -2708 -7676 -2702
rect -7718 -2727 -7715 -2712
rect -7684 -2712 -7676 -2708
rect -7707 -2720 -7692 -2716
rect -7723 -2773 -7714 -2769
rect -7704 -2770 -7700 -2720
rect -7680 -2727 -7676 -2712
rect -7583 -2714 -7580 -2708
rect -7583 -2718 -7576 -2714
rect -7569 -2715 -7565 -2684
rect -7545 -2714 -7541 -2708
rect -7583 -2733 -7580 -2718
rect -7549 -2718 -7541 -2714
rect -7572 -2726 -7557 -2722
rect -7957 -2803 -7949 -2799
rect -7942 -2800 -7938 -2790
rect -7864 -2798 -7860 -2789
rect -7857 -2797 -7853 -2780
rect -7815 -2780 -7807 -2776
rect -7844 -2788 -7823 -2784
rect -7857 -2801 -7848 -2797
rect -7957 -2811 -7949 -2807
rect -7953 -2820 -7949 -2811
rect -7857 -2809 -7848 -2805
rect -7857 -2818 -7853 -2809
rect -7956 -2848 -7952 -2842
rect -7994 -2867 -7991 -2852
rect -7960 -2852 -7952 -2848
rect -7983 -2860 -7968 -2856
rect -8126 -2892 -8110 -2888
rect -8087 -2889 -8083 -2877
rect -8002 -2892 -7998 -2878
rect -7980 -2891 -7976 -2860
rect -7956 -2867 -7952 -2852
rect -7852 -2846 -7849 -2840
rect -7852 -2850 -7845 -2846
rect -7838 -2847 -7834 -2788
rect -7811 -2797 -7807 -2780
rect -7815 -2801 -7807 -2797
rect -7800 -2798 -7796 -2788
rect -7730 -2791 -7726 -2782
rect -7723 -2790 -7719 -2773
rect -7681 -2773 -7673 -2769
rect -7710 -2781 -7689 -2777
rect -7723 -2794 -7714 -2790
rect -7723 -2802 -7714 -2798
rect -7815 -2809 -7807 -2805
rect -7811 -2818 -7807 -2809
rect -7723 -2811 -7719 -2802
rect -7718 -2839 -7715 -2833
rect -7814 -2846 -7810 -2840
rect -7852 -2865 -7849 -2850
rect -7818 -2850 -7810 -2846
rect -7841 -2858 -7826 -2854
rect -7984 -2895 -7968 -2891
rect -7945 -2892 -7941 -2880
rect -7860 -2890 -7856 -2876
rect -7838 -2889 -7834 -2858
rect -7814 -2865 -7810 -2850
rect -7718 -2843 -7711 -2839
rect -7704 -2840 -7700 -2781
rect -7677 -2790 -7673 -2773
rect -7588 -2779 -7579 -2775
rect -7569 -2776 -7565 -2726
rect -7545 -2733 -7541 -2718
rect -7463 -2713 -7460 -2707
rect -7463 -2717 -7456 -2713
rect -7449 -2714 -7445 -2683
rect -7425 -2713 -7421 -2707
rect -7463 -2732 -7460 -2717
rect -7429 -2717 -7421 -2713
rect -7452 -2725 -7437 -2721
rect -7681 -2794 -7673 -2790
rect -7666 -2791 -7662 -2781
rect -7595 -2797 -7591 -2788
rect -7681 -2802 -7673 -2798
rect -7588 -2796 -7584 -2779
rect -7546 -2779 -7538 -2775
rect -7575 -2787 -7554 -2783
rect -7588 -2800 -7579 -2796
rect -7677 -2811 -7673 -2802
rect -7588 -2808 -7579 -2804
rect -7588 -2817 -7584 -2808
rect -7680 -2839 -7676 -2833
rect -7718 -2858 -7715 -2843
rect -7684 -2843 -7676 -2839
rect -7707 -2851 -7692 -2847
rect -7842 -2893 -7826 -2889
rect -7803 -2890 -7799 -2878
rect -7726 -2883 -7722 -2869
rect -7704 -2882 -7700 -2851
rect -7680 -2858 -7676 -2843
rect -7583 -2845 -7580 -2839
rect -7583 -2849 -7576 -2845
rect -7569 -2846 -7565 -2787
rect -7542 -2796 -7538 -2779
rect -7468 -2778 -7459 -2774
rect -7449 -2775 -7445 -2725
rect -7425 -2732 -7421 -2717
rect -7343 -2713 -7340 -2707
rect -7343 -2717 -7336 -2713
rect -7329 -2714 -7325 -2683
rect -7305 -2713 -7301 -2707
rect -7343 -2732 -7340 -2717
rect -7309 -2717 -7301 -2713
rect -7332 -2725 -7317 -2721
rect -7546 -2800 -7538 -2796
rect -7531 -2797 -7527 -2787
rect -7475 -2796 -7471 -2787
rect -7468 -2795 -7464 -2778
rect -7426 -2778 -7418 -2774
rect -7455 -2786 -7434 -2782
rect -7468 -2799 -7459 -2795
rect -7546 -2808 -7538 -2804
rect -7542 -2817 -7538 -2808
rect -7468 -2807 -7459 -2803
rect -7468 -2816 -7464 -2807
rect -7545 -2845 -7541 -2839
rect -7583 -2864 -7580 -2849
rect -7549 -2849 -7541 -2845
rect -7572 -2857 -7557 -2853
rect -7708 -2886 -7692 -2882
rect -7669 -2883 -7665 -2871
rect -7591 -2889 -7587 -2875
rect -7569 -2888 -7565 -2857
rect -7545 -2864 -7541 -2849
rect -7463 -2844 -7460 -2838
rect -7463 -2848 -7456 -2844
rect -7449 -2845 -7445 -2786
rect -7422 -2795 -7418 -2778
rect -7348 -2778 -7339 -2774
rect -7329 -2775 -7325 -2725
rect -7305 -2732 -7301 -2717
rect -7218 -2712 -7215 -2706
rect -7218 -2716 -7211 -2712
rect -7204 -2713 -7200 -2682
rect -7180 -2712 -7176 -2706
rect -7218 -2731 -7215 -2716
rect -7184 -2716 -7176 -2712
rect -7207 -2724 -7192 -2720
rect -7426 -2799 -7418 -2795
rect -7411 -2796 -7407 -2786
rect -7355 -2796 -7351 -2787
rect -7348 -2795 -7344 -2778
rect -7306 -2778 -7298 -2774
rect -7335 -2786 -7314 -2782
rect -7348 -2799 -7339 -2795
rect -7426 -2807 -7418 -2803
rect -7422 -2816 -7418 -2807
rect -7348 -2807 -7339 -2803
rect -7348 -2816 -7344 -2807
rect -7425 -2844 -7421 -2838
rect -7463 -2863 -7460 -2848
rect -7429 -2848 -7421 -2844
rect -7452 -2856 -7437 -2852
rect -7708 -2894 -7692 -2890
rect -7573 -2892 -7557 -2888
rect -7534 -2889 -7530 -2877
rect -7471 -2888 -7467 -2874
rect -7449 -2887 -7445 -2856
rect -7425 -2863 -7421 -2848
rect -7343 -2844 -7340 -2838
rect -7343 -2848 -7336 -2844
rect -7329 -2845 -7325 -2786
rect -7302 -2795 -7298 -2778
rect -7223 -2777 -7214 -2773
rect -7204 -2774 -7200 -2724
rect -7180 -2731 -7176 -2716
rect -7100 -2712 -7097 -2706
rect -7100 -2716 -7093 -2712
rect -7086 -2713 -7082 -2682
rect -7062 -2712 -7058 -2706
rect -7100 -2731 -7097 -2716
rect -7066 -2716 -7058 -2712
rect -7089 -2724 -7074 -2720
rect -7306 -2799 -7298 -2795
rect -7291 -2796 -7287 -2786
rect -7230 -2795 -7226 -2786
rect -7223 -2794 -7219 -2777
rect -7181 -2777 -7173 -2773
rect -7210 -2785 -7189 -2781
rect -7223 -2798 -7214 -2794
rect -7306 -2807 -7298 -2803
rect -7302 -2816 -7298 -2807
rect -7223 -2806 -7214 -2802
rect -7223 -2815 -7219 -2806
rect -7305 -2844 -7301 -2838
rect -7343 -2863 -7340 -2848
rect -7309 -2848 -7301 -2844
rect -7332 -2856 -7317 -2852
rect -7453 -2891 -7437 -2887
rect -7414 -2888 -7410 -2876
rect -7351 -2888 -7347 -2874
rect -7329 -2887 -7325 -2856
rect -7305 -2863 -7301 -2848
rect -7218 -2843 -7215 -2837
rect -7218 -2847 -7211 -2843
rect -7204 -2844 -7200 -2785
rect -7177 -2794 -7173 -2777
rect -7105 -2777 -7096 -2773
rect -7086 -2774 -7082 -2724
rect -7062 -2731 -7058 -2716
rect -6981 -2710 -6978 -2704
rect -6981 -2714 -6974 -2710
rect -6967 -2711 -6963 -2680
rect -6943 -2710 -6939 -2704
rect -6981 -2729 -6978 -2714
rect -6947 -2714 -6939 -2710
rect -6970 -2722 -6955 -2718
rect -7181 -2798 -7173 -2794
rect -7166 -2795 -7162 -2785
rect -7112 -2795 -7108 -2786
rect -7105 -2794 -7101 -2777
rect -7063 -2777 -7055 -2773
rect -7092 -2785 -7071 -2781
rect -7105 -2798 -7096 -2794
rect -7181 -2806 -7173 -2802
rect -7177 -2815 -7173 -2806
rect -7105 -2806 -7096 -2802
rect -7105 -2815 -7101 -2806
rect -7180 -2843 -7176 -2837
rect -7218 -2862 -7215 -2847
rect -7184 -2847 -7176 -2843
rect -7207 -2855 -7192 -2851
rect -7333 -2891 -7317 -2887
rect -7294 -2888 -7290 -2876
rect -7226 -2887 -7222 -2873
rect -7204 -2886 -7200 -2855
rect -7180 -2862 -7176 -2847
rect -7100 -2843 -7097 -2837
rect -7100 -2847 -7093 -2843
rect -7086 -2844 -7082 -2785
rect -7059 -2794 -7055 -2777
rect -6986 -2775 -6977 -2771
rect -6967 -2772 -6963 -2722
rect -6943 -2729 -6939 -2714
rect -7063 -2798 -7055 -2794
rect -7048 -2795 -7044 -2785
rect -6993 -2793 -6989 -2784
rect -6986 -2792 -6982 -2775
rect -6944 -2775 -6936 -2771
rect -6973 -2783 -6952 -2779
rect -6986 -2796 -6977 -2792
rect -7063 -2806 -7055 -2802
rect -7059 -2815 -7055 -2806
rect -6986 -2804 -6977 -2800
rect -6986 -2813 -6982 -2804
rect -7062 -2843 -7058 -2837
rect -7100 -2862 -7097 -2847
rect -7066 -2847 -7058 -2843
rect -7089 -2855 -7074 -2851
rect -7208 -2890 -7192 -2886
rect -7169 -2887 -7165 -2875
rect -7108 -2887 -7104 -2873
rect -7086 -2886 -7082 -2855
rect -7062 -2862 -7058 -2847
rect -6981 -2841 -6978 -2835
rect -6981 -2845 -6974 -2841
rect -6967 -2842 -6963 -2783
rect -6940 -2792 -6936 -2775
rect -6944 -2796 -6936 -2792
rect -6929 -2793 -6925 -2783
rect -6944 -2804 -6936 -2800
rect -6940 -2813 -6936 -2804
rect -6943 -2841 -6939 -2835
rect -6981 -2860 -6978 -2845
rect -6947 -2845 -6939 -2841
rect -6970 -2853 -6955 -2849
rect -7090 -2890 -7074 -2886
rect -7051 -2887 -7047 -2875
rect -6989 -2885 -6985 -2871
rect -6967 -2884 -6963 -2853
rect -6943 -2860 -6939 -2845
rect -6971 -2888 -6955 -2884
rect -6932 -2885 -6928 -2873
rect -8126 -2900 -8110 -2896
rect -8136 -2930 -8133 -2924
rect -8136 -2934 -8129 -2930
rect -8122 -2931 -8118 -2900
rect -7984 -2903 -7968 -2899
rect -7842 -2901 -7826 -2897
rect -8098 -2930 -8094 -2924
rect -8136 -2949 -8133 -2934
rect -8102 -2934 -8094 -2930
rect -8125 -2942 -8110 -2938
rect -8141 -2995 -8132 -2991
rect -8122 -2992 -8118 -2942
rect -8098 -2949 -8094 -2934
rect -7994 -2933 -7991 -2927
rect -7994 -2937 -7987 -2933
rect -7980 -2934 -7976 -2903
rect -7956 -2933 -7952 -2927
rect -7994 -2952 -7991 -2937
rect -7960 -2937 -7952 -2933
rect -7983 -2945 -7968 -2941
rect -8148 -3013 -8144 -3004
rect -8141 -3012 -8137 -2995
rect -8099 -2995 -8091 -2991
rect -8128 -3003 -8107 -2999
rect -8141 -3016 -8132 -3012
rect -8141 -3024 -8132 -3020
rect -8141 -3033 -8137 -3024
rect -8122 -3043 -8118 -3003
rect -8095 -3012 -8091 -2995
rect -7999 -2998 -7990 -2994
rect -7980 -2995 -7976 -2945
rect -7956 -2952 -7952 -2937
rect -7852 -2931 -7849 -2925
rect -7852 -2935 -7845 -2931
rect -7838 -2932 -7834 -2901
rect -7718 -2924 -7715 -2918
rect -7814 -2931 -7810 -2925
rect -7852 -2950 -7849 -2935
rect -7818 -2935 -7810 -2931
rect -7841 -2943 -7826 -2939
rect -8099 -3016 -8091 -3012
rect -8084 -3013 -8080 -3003
rect -8006 -3016 -8002 -3007
rect -7999 -3015 -7995 -2998
rect -7957 -2998 -7949 -2994
rect -7986 -3006 -7965 -3002
rect -7999 -3019 -7990 -3015
rect -8099 -3024 -8091 -3020
rect -8095 -3033 -8091 -3024
rect -7999 -3027 -7990 -3023
rect -7999 -3036 -7995 -3027
rect -7980 -3049 -7976 -3006
rect -7953 -3015 -7949 -2998
rect -7857 -2996 -7848 -2992
rect -7838 -2993 -7834 -2943
rect -7814 -2950 -7810 -2935
rect -7718 -2928 -7711 -2924
rect -7704 -2925 -7700 -2894
rect -7573 -2900 -7557 -2896
rect -7453 -2899 -7437 -2895
rect -7333 -2899 -7317 -2895
rect -7208 -2898 -7192 -2894
rect -7090 -2898 -7074 -2894
rect -6971 -2896 -6955 -2892
rect -7680 -2924 -7676 -2918
rect -7718 -2943 -7715 -2928
rect -7684 -2928 -7676 -2924
rect -7707 -2936 -7692 -2932
rect -7723 -2989 -7714 -2985
rect -7704 -2986 -7700 -2936
rect -7680 -2943 -7676 -2928
rect -7583 -2930 -7580 -2924
rect -7583 -2934 -7576 -2930
rect -7569 -2931 -7565 -2900
rect -7545 -2930 -7541 -2924
rect -7583 -2949 -7580 -2934
rect -7549 -2934 -7541 -2930
rect -7572 -2942 -7557 -2938
rect -7957 -3019 -7949 -3015
rect -7942 -3016 -7938 -3006
rect -7864 -3014 -7860 -3005
rect -7857 -3013 -7853 -2996
rect -7815 -2996 -7807 -2992
rect -7844 -3004 -7823 -3000
rect -7857 -3017 -7848 -3013
rect -7957 -3027 -7949 -3023
rect -7953 -3036 -7949 -3027
rect -7857 -3025 -7848 -3021
rect -7857 -3034 -7853 -3025
rect -7838 -3047 -7834 -3004
rect -7811 -3013 -7807 -2996
rect -7815 -3017 -7807 -3013
rect -7800 -3014 -7796 -3004
rect -7730 -3007 -7726 -2998
rect -7723 -3006 -7719 -2989
rect -7681 -2989 -7673 -2985
rect -7710 -2997 -7689 -2993
rect -7723 -3010 -7714 -3006
rect -7723 -3018 -7714 -3014
rect -7815 -3025 -7807 -3021
rect -7811 -3034 -7807 -3025
rect -7723 -3027 -7719 -3018
rect -7704 -3036 -7700 -2997
rect -7677 -3006 -7673 -2989
rect -7588 -2995 -7579 -2991
rect -7569 -2992 -7565 -2942
rect -7545 -2949 -7541 -2934
rect -7463 -2929 -7460 -2923
rect -7463 -2933 -7456 -2929
rect -7449 -2930 -7445 -2899
rect -7425 -2929 -7421 -2923
rect -7463 -2948 -7460 -2933
rect -7429 -2933 -7421 -2929
rect -7452 -2941 -7437 -2937
rect -7681 -3010 -7673 -3006
rect -7666 -3007 -7662 -2997
rect -7595 -3013 -7591 -3004
rect -7681 -3018 -7673 -3014
rect -7588 -3012 -7584 -2995
rect -7546 -2995 -7538 -2991
rect -7575 -3003 -7554 -2999
rect -7588 -3016 -7579 -3012
rect -7677 -3027 -7673 -3018
rect -7588 -3024 -7579 -3020
rect -7588 -3033 -7584 -3024
rect -7569 -3046 -7565 -3003
rect -7542 -3012 -7538 -2995
rect -7468 -2994 -7459 -2990
rect -7449 -2991 -7445 -2941
rect -7425 -2948 -7421 -2933
rect -7343 -2929 -7340 -2923
rect -7343 -2933 -7336 -2929
rect -7329 -2930 -7325 -2899
rect -7305 -2929 -7301 -2923
rect -7343 -2948 -7340 -2933
rect -7309 -2933 -7301 -2929
rect -7332 -2941 -7317 -2937
rect -7546 -3016 -7538 -3012
rect -7531 -3013 -7527 -3003
rect -7475 -3012 -7471 -3003
rect -7468 -3011 -7464 -2994
rect -7426 -2994 -7418 -2990
rect -7455 -3002 -7434 -2998
rect -7468 -3015 -7459 -3011
rect -7546 -3024 -7538 -3020
rect -7542 -3033 -7538 -3024
rect -7468 -3023 -7459 -3019
rect -7468 -3032 -7464 -3023
rect -7449 -3038 -7445 -3002
rect -7422 -3011 -7418 -2994
rect -7348 -2994 -7339 -2990
rect -7329 -2991 -7325 -2941
rect -7305 -2948 -7301 -2933
rect -7218 -2928 -7215 -2922
rect -7218 -2932 -7211 -2928
rect -7204 -2929 -7200 -2898
rect -7180 -2928 -7176 -2922
rect -7218 -2947 -7215 -2932
rect -7184 -2932 -7176 -2928
rect -7207 -2940 -7192 -2936
rect -7426 -3015 -7418 -3011
rect -7411 -3012 -7407 -3002
rect -7355 -3012 -7351 -3003
rect -7348 -3011 -7344 -2994
rect -7306 -2994 -7298 -2990
rect -7335 -3002 -7314 -2998
rect -7348 -3015 -7339 -3011
rect -7426 -3023 -7418 -3019
rect -7422 -3032 -7418 -3023
rect -7348 -3023 -7339 -3019
rect -7348 -3032 -7344 -3023
rect -7329 -3038 -7325 -3002
rect -7302 -3011 -7298 -2994
rect -7223 -2993 -7214 -2989
rect -7204 -2990 -7200 -2940
rect -7180 -2947 -7176 -2932
rect -7100 -2928 -7097 -2922
rect -7100 -2932 -7093 -2928
rect -7086 -2929 -7082 -2898
rect -7062 -2928 -7058 -2922
rect -7100 -2947 -7097 -2932
rect -7066 -2932 -7058 -2928
rect -7089 -2940 -7074 -2936
rect -7306 -3015 -7298 -3011
rect -7291 -3012 -7287 -3002
rect -7230 -3011 -7226 -3002
rect -7223 -3010 -7219 -2993
rect -7181 -2993 -7173 -2989
rect -7210 -3001 -7189 -2997
rect -7223 -3014 -7214 -3010
rect -7306 -3023 -7298 -3019
rect -7302 -3032 -7298 -3023
rect -7223 -3022 -7214 -3018
rect -7223 -3031 -7219 -3022
rect -7204 -3037 -7200 -3001
rect -7177 -3010 -7173 -2993
rect -7105 -2993 -7096 -2989
rect -7086 -2990 -7082 -2940
rect -7062 -2947 -7058 -2932
rect -6981 -2926 -6978 -2920
rect -6981 -2930 -6974 -2926
rect -6967 -2927 -6963 -2896
rect -6943 -2926 -6939 -2920
rect -6981 -2945 -6978 -2930
rect -6947 -2930 -6939 -2926
rect -6970 -2938 -6955 -2934
rect -7181 -3014 -7173 -3010
rect -7166 -3011 -7162 -3001
rect -7112 -3011 -7108 -3002
rect -7105 -3010 -7101 -2993
rect -7063 -2993 -7055 -2989
rect -7092 -3001 -7071 -2997
rect -7105 -3014 -7096 -3010
rect -7181 -3022 -7173 -3018
rect -7177 -3031 -7173 -3022
rect -7105 -3022 -7096 -3018
rect -7105 -3031 -7101 -3022
rect -7086 -3037 -7082 -3001
rect -7059 -3010 -7055 -2993
rect -6986 -2991 -6977 -2987
rect -6967 -2988 -6963 -2938
rect -6943 -2945 -6939 -2930
rect -7063 -3014 -7055 -3010
rect -7048 -3011 -7044 -3001
rect -6993 -3009 -6989 -3000
rect -6986 -3008 -6982 -2991
rect -6944 -2991 -6936 -2987
rect -6973 -2999 -6952 -2995
rect -6986 -3012 -6977 -3008
rect -7063 -3022 -7055 -3018
rect -7059 -3031 -7055 -3022
rect -6986 -3020 -6977 -3016
rect -6986 -3029 -6982 -3020
rect -6967 -3035 -6963 -2999
rect -6940 -3008 -6936 -2991
rect -6944 -3012 -6936 -3008
rect -6929 -3009 -6925 -2999
rect -6944 -3020 -6936 -3016
rect -6940 -3029 -6936 -3020
rect -7449 -3050 -7446 -3038
rect -7329 -3050 -7326 -3038
rect -7449 -4153 -7445 -3050
rect -7329 -3937 -7325 -3050
rect -7204 -3789 -7201 -3037
rect -7086 -3048 -7083 -3037
rect -7086 -3645 -7082 -3048
rect -6967 -3473 -6964 -3035
rect -5882 -3169 -5877 -2602
rect -6316 -3174 -5877 -3169
rect -6078 -3446 -6050 -3443
rect -6077 -3452 -6074 -3446
rect -6053 -3447 -6050 -3446
rect -6053 -3450 -5982 -3447
rect -6373 -3473 -6368 -3472
rect -6967 -3476 -6091 -3473
rect -6373 -3477 -6368 -3476
rect -6086 -3475 -6076 -3472
rect -6068 -3472 -6065 -3464
rect -6038 -3456 -6035 -3450
rect -6019 -3456 -6016 -3450
rect -6068 -3475 -6047 -3472
rect -6068 -3478 -6065 -3475
rect -6077 -3488 -6074 -3484
rect -6083 -3490 -6059 -3488
rect -6083 -3491 -6065 -3490
rect -6060 -3491 -6059 -3490
rect -6050 -3498 -6047 -3475
rect -6009 -3456 -5989 -3453
rect -6009 -3462 -6006 -3456
rect -5992 -3462 -5989 -3456
rect -6028 -3483 -6025 -3480
rect -6028 -3486 -6010 -3483
rect -6000 -3493 -5997 -3486
rect -6000 -3496 -5983 -3493
rect -6078 -3499 -6059 -3498
rect -6083 -3501 -6059 -3499
rect -6050 -3501 -6007 -3498
rect -6077 -3507 -6074 -3501
rect -5986 -3507 -5983 -3496
rect -6021 -3512 -5996 -3509
rect -5986 -3510 -5972 -3507
rect -5986 -3511 -5977 -3510
rect -6021 -3514 -6018 -3512
rect -6271 -3530 -6091 -3527
rect -6086 -3530 -6076 -3527
rect -6068 -3527 -6065 -3519
rect -6056 -3517 -6018 -3514
rect -5986 -3515 -5983 -3511
rect -6056 -3527 -6053 -3517
rect -6015 -3518 -5983 -3515
rect -6015 -3521 -6012 -3518
rect -6068 -3530 -6053 -3527
rect -6068 -3533 -6065 -3530
rect -6016 -3524 -6010 -3521
rect -6077 -3543 -6074 -3539
rect -6056 -3540 -6051 -3537
rect -6038 -3537 -6035 -3533
rect -5991 -3537 -5988 -3533
rect -6046 -3540 -5982 -3537
rect -6056 -3543 -6053 -3540
rect -6083 -3546 -6053 -3543
rect -6085 -3618 -6057 -3615
rect -6084 -3624 -6081 -3618
rect -6060 -3619 -6057 -3618
rect -6060 -3622 -5989 -3619
rect -7086 -3648 -6098 -3645
rect -7086 -3650 -6180 -3648
rect -6093 -3647 -6083 -3644
rect -6075 -3644 -6072 -3636
rect -6045 -3628 -6042 -3622
rect -6026 -3628 -6023 -3622
rect -6075 -3647 -6054 -3644
rect -6075 -3650 -6072 -3647
rect -6084 -3660 -6081 -3656
rect -6090 -3662 -6066 -3660
rect -6090 -3663 -6072 -3662
rect -6067 -3663 -6066 -3662
rect -6057 -3670 -6054 -3647
rect -6016 -3628 -5996 -3625
rect -6016 -3634 -6013 -3628
rect -5999 -3634 -5996 -3628
rect -6035 -3655 -6032 -3652
rect -6035 -3658 -6017 -3655
rect -6007 -3665 -6004 -3658
rect -6007 -3668 -5990 -3665
rect -6085 -3671 -6066 -3670
rect -6090 -3673 -6066 -3671
rect -6057 -3673 -6014 -3670
rect -6084 -3679 -6081 -3673
rect -5993 -3679 -5990 -3668
rect -5984 -3679 -5979 -3604
rect -6028 -3684 -6003 -3681
rect -5993 -3683 -5979 -3679
rect -6028 -3686 -6025 -3684
rect -6180 -3702 -6098 -3699
rect -6093 -3702 -6083 -3699
rect -6075 -3699 -6072 -3691
rect -6063 -3689 -6025 -3686
rect -5993 -3687 -5990 -3683
rect -6063 -3699 -6060 -3689
rect -6022 -3690 -5990 -3687
rect -6022 -3693 -6019 -3690
rect -6075 -3702 -6060 -3699
rect -6075 -3705 -6072 -3702
rect -6023 -3696 -6017 -3693
rect -6084 -3715 -6081 -3711
rect -6063 -3712 -6058 -3709
rect -6045 -3709 -6042 -3705
rect -5998 -3709 -5995 -3705
rect -6053 -3712 -5989 -3709
rect -6063 -3715 -6060 -3712
rect -6090 -3718 -6060 -3715
rect -6082 -3762 -6054 -3759
rect -6081 -3768 -6078 -3762
rect -6057 -3763 -6054 -3762
rect -6057 -3766 -5986 -3763
rect -7204 -3792 -6095 -3789
rect -7204 -3794 -6170 -3792
rect -6090 -3791 -6080 -3788
rect -6072 -3788 -6069 -3780
rect -6042 -3772 -6039 -3766
rect -6023 -3772 -6020 -3766
rect -6072 -3791 -6051 -3788
rect -6072 -3794 -6069 -3791
rect -6081 -3804 -6078 -3800
rect -6087 -3806 -6063 -3804
rect -6087 -3807 -6069 -3806
rect -6064 -3807 -6063 -3806
rect -6054 -3814 -6051 -3791
rect -6013 -3772 -5993 -3769
rect -6013 -3778 -6010 -3772
rect -5996 -3778 -5993 -3772
rect -5882 -3778 -5877 -3174
rect -5765 -3510 -5760 -2666
rect -5708 -3599 -5703 -2752
rect -6032 -3799 -6029 -3796
rect -6032 -3802 -6014 -3799
rect -6004 -3809 -6001 -3802
rect -6004 -3812 -5987 -3809
rect -6082 -3815 -6063 -3814
rect -6087 -3817 -6063 -3815
rect -6054 -3817 -6011 -3814
rect -6081 -3823 -6078 -3817
rect -5990 -3823 -5987 -3812
rect -6025 -3828 -6000 -3825
rect -5990 -3827 -5976 -3823
rect -6025 -3830 -6022 -3828
rect -6178 -3846 -6095 -3843
rect -6090 -3846 -6080 -3843
rect -6072 -3843 -6069 -3835
rect -6060 -3833 -6022 -3830
rect -5990 -3831 -5987 -3827
rect -6060 -3843 -6057 -3833
rect -6019 -3834 -5987 -3831
rect -5981 -3833 -5976 -3827
rect -6019 -3837 -6016 -3834
rect -6072 -3846 -6057 -3843
rect -6072 -3849 -6069 -3846
rect -6020 -3840 -6014 -3837
rect -5616 -3833 -5611 -2813
rect -6081 -3859 -6078 -3855
rect -6060 -3856 -6055 -3853
rect -6042 -3853 -6039 -3849
rect -5995 -3853 -5992 -3849
rect -6050 -3856 -5986 -3853
rect -6060 -3859 -6057 -3856
rect -6087 -3862 -6057 -3859
rect -5487 -3864 -5482 -2902
rect -6086 -3910 -6058 -3907
rect -6085 -3916 -6082 -3910
rect -6061 -3911 -6058 -3910
rect -6061 -3914 -5990 -3911
rect -7329 -3940 -6099 -3937
rect -7329 -3942 -6172 -3940
rect -6094 -3939 -6084 -3936
rect -6076 -3936 -6073 -3928
rect -6046 -3920 -6043 -3914
rect -6027 -3920 -6024 -3914
rect -6076 -3939 -6055 -3936
rect -6076 -3942 -6073 -3939
rect -6085 -3952 -6082 -3948
rect -6091 -3954 -6067 -3952
rect -6091 -3955 -6073 -3954
rect -6068 -3955 -6067 -3954
rect -6058 -3962 -6055 -3939
rect -6017 -3920 -5997 -3917
rect -6017 -3926 -6014 -3920
rect -6000 -3926 -5997 -3920
rect -6036 -3947 -6033 -3944
rect -6036 -3950 -6018 -3947
rect -6008 -3957 -6005 -3950
rect -6008 -3960 -5991 -3957
rect -6086 -3963 -6067 -3962
rect -6091 -3965 -6067 -3963
rect -6058 -3965 -6015 -3962
rect -6085 -3971 -6082 -3965
rect -5994 -3971 -5991 -3960
rect -5985 -3971 -5980 -3869
rect -6029 -3976 -6004 -3973
rect -5994 -3975 -5980 -3971
rect -6029 -3978 -6026 -3976
rect -6174 -3994 -6099 -3991
rect -6094 -3994 -6084 -3991
rect -6076 -3991 -6073 -3983
rect -6064 -3981 -6026 -3978
rect -5994 -3979 -5991 -3975
rect -6064 -3991 -6061 -3981
rect -6023 -3982 -5991 -3979
rect -6023 -3985 -6020 -3982
rect -6076 -3994 -6061 -3991
rect -6076 -3997 -6073 -3994
rect -6024 -3988 -6018 -3985
rect -6085 -4007 -6082 -4003
rect -6064 -4004 -6059 -4001
rect -6046 -4001 -6043 -3997
rect -5999 -4001 -5996 -3997
rect -6054 -4004 -5990 -4001
rect -6064 -4007 -6061 -4004
rect -6091 -4010 -6061 -4007
rect -5327 -4027 -5322 -2947
rect -5237 -2980 -5233 -2977
rect -5243 -2984 -5242 -2980
rect -5238 -2984 -5233 -2980
rect -5237 -2990 -5233 -2984
rect -5229 -3040 -5225 -3030
rect -5229 -3046 -5189 -3040
rect -5229 -3048 -5225 -3046
rect -5237 -3078 -5233 -3068
rect -5196 -3151 -5189 -3046
rect -5196 -3154 -4684 -3151
rect -5196 -3157 -4544 -3154
rect -5196 -3284 -5189 -3157
rect -5103 -3206 -5099 -3197
rect -5109 -3211 -5108 -3206
rect -5104 -3211 -5085 -3206
rect -5103 -3217 -5099 -3211
rect -5196 -3290 -5115 -3284
rect -5196 -3292 -5189 -3290
rect -5095 -3320 -5091 -3267
rect -4981 -3285 -4974 -3157
rect -4931 -3207 -4927 -3198
rect -4937 -3212 -4936 -3207
rect -4932 -3212 -4913 -3207
rect -4931 -3218 -4927 -3212
rect -4981 -3291 -4942 -3285
rect -5095 -3325 -4992 -3320
rect -5095 -3399 -5091 -3325
rect -4997 -3399 -4992 -3325
rect -5087 -3667 -5083 -3499
rect -4997 -3637 -4992 -3404
rect -4923 -3327 -4919 -3268
rect -4811 -3285 -4805 -3157
rect -4690 -3160 -4544 -3157
rect -4757 -3207 -4753 -3198
rect -4763 -3212 -4762 -3207
rect -4758 -3212 -4739 -3207
rect -4757 -3218 -4753 -3212
rect -4811 -3291 -4768 -3285
rect -4749 -3322 -4745 -3268
rect -4690 -3286 -4684 -3160
rect -4633 -3208 -4629 -3199
rect -4639 -3213 -4638 -3208
rect -4634 -3213 -4615 -3208
rect -4633 -3219 -4629 -3213
rect -4690 -3292 -4644 -3286
rect -4749 -3327 -4652 -3322
rect -4923 -3332 -4809 -3327
rect -4923 -3488 -4919 -3332
rect -4915 -3637 -4911 -3588
rect -4997 -3644 -4911 -3637
rect -6061 -4126 -6033 -4123
rect -6060 -4132 -6057 -4126
rect -6036 -4127 -6033 -4126
rect -6036 -4130 -5965 -4127
rect -7449 -4156 -6074 -4153
rect -7449 -4158 -6149 -4156
rect -6069 -4155 -6059 -4152
rect -6051 -4152 -6048 -4144
rect -6021 -4136 -6018 -4130
rect -6002 -4136 -5999 -4130
rect -6051 -4155 -6030 -4152
rect -6051 -4158 -6048 -4155
rect -6060 -4168 -6057 -4164
rect -6066 -4170 -6042 -4168
rect -6066 -4171 -6048 -4170
rect -6043 -4171 -6042 -4170
rect -6033 -4178 -6030 -4155
rect -5992 -4136 -5972 -4133
rect -5992 -4142 -5989 -4136
rect -5975 -4142 -5972 -4136
rect -6011 -4163 -6008 -4160
rect -6011 -4166 -5993 -4163
rect -5983 -4173 -5980 -4166
rect -5983 -4176 -5966 -4173
rect -6061 -4179 -6042 -4178
rect -6066 -4181 -6042 -4179
rect -6033 -4181 -5990 -4178
rect -6060 -4187 -6057 -4181
rect -5969 -4187 -5966 -4176
rect -5960 -4187 -5955 -4032
rect -6004 -4192 -5979 -4189
rect -5969 -4191 -5955 -4187
rect -6004 -4194 -6001 -4192
rect -6149 -4210 -6074 -4207
rect -6069 -4210 -6059 -4207
rect -6051 -4207 -6048 -4199
rect -6039 -4197 -6001 -4194
rect -5969 -4195 -5966 -4191
rect -6039 -4207 -6036 -4197
rect -5998 -4198 -5966 -4195
rect -5998 -4201 -5995 -4198
rect -6051 -4210 -6036 -4207
rect -6051 -4213 -6048 -4210
rect -5999 -4204 -5993 -4201
rect -6060 -4223 -6057 -4219
rect -6039 -4220 -6034 -4217
rect -6021 -4217 -6018 -4213
rect -5974 -4217 -5971 -4213
rect -6029 -4220 -5965 -4217
rect -6039 -4223 -6036 -4220
rect -6066 -4226 -6036 -4223
rect -5079 -4269 -5075 -3767
rect -4915 -4269 -4911 -3644
rect -4814 -3530 -4809 -3332
rect -4814 -3891 -4809 -3535
rect -4749 -3722 -4745 -3327
rect -4657 -3661 -4652 -3327
rect -4741 -3891 -4737 -3822
rect -4814 -3896 -4737 -3891
rect -4741 -4269 -4737 -3896
rect -4657 -3903 -4652 -3666
rect -4625 -3359 -4621 -3269
rect -4550 -3289 -4544 -3160
rect -4493 -3211 -4489 -3202
rect -4499 -3216 -4498 -3211
rect -4494 -3216 -4475 -3211
rect -4493 -3222 -4489 -3216
rect -4550 -3295 -4504 -3289
rect -4485 -3359 -4481 -3272
rect -4294 -3339 -4290 -3336
rect -4300 -3343 -4299 -3339
rect -4295 -3343 -4290 -3339
rect -4294 -3349 -4290 -3343
rect -4625 -3364 -4535 -3359
rect -4625 -3753 -4621 -3364
rect -4617 -3903 -4613 -3853
rect -4657 -3908 -4613 -3903
rect -4617 -4269 -4613 -3908
rect -4540 -3804 -4535 -3364
rect -4540 -4046 -4535 -3809
rect -4485 -3365 -4393 -3359
rect -4485 -3916 -4481 -3365
rect -4477 -4046 -4473 -4016
rect -4540 -4050 -4473 -4046
rect -6061 -4364 -6038 -4360
rect -6057 -4366 -6038 -4364
rect -6061 -4375 -6057 -4370
rect -6042 -4375 -6038 -4366
rect -6025 -4371 -6001 -4370
rect -6025 -4375 -6009 -4371
rect -6005 -4375 -6001 -4371
rect -6025 -4377 -6001 -4375
rect -6019 -4382 -6015 -4377
rect -6050 -4403 -6046 -4395
rect -6050 -4407 -6038 -4403
rect -6042 -4409 -6038 -4407
rect -6011 -4409 -6007 -4402
rect -5990 -4409 -5984 -4407
rect -6208 -4414 -6049 -4410
rect -6042 -4413 -6018 -4409
rect -6011 -4413 -5984 -4409
rect -6219 -4418 -6060 -4417
rect -6213 -4421 -6060 -4418
rect -6042 -4424 -6038 -4413
rect -6011 -4416 -6007 -4413
rect -6019 -4430 -6015 -4426
rect -6025 -4431 -6000 -4430
rect -6025 -4435 -6005 -4431
rect -6025 -4436 -6000 -4435
rect -6061 -4448 -6057 -4444
rect -6061 -4452 -6045 -4448
rect -6060 -4473 -6037 -4469
rect -6056 -4475 -6037 -4473
rect -6060 -4484 -6056 -4479
rect -6041 -4484 -6037 -4475
rect -6024 -4480 -6000 -4479
rect -6024 -4484 -6008 -4480
rect -6004 -4484 -6000 -4480
rect -6024 -4486 -6000 -4484
rect -6018 -4491 -6014 -4486
rect -6049 -4512 -6045 -4504
rect -6049 -4516 -6037 -4512
rect -6041 -4518 -6037 -4516
rect -6010 -4518 -6006 -4511
rect -5996 -4518 -5991 -4440
rect -6115 -4523 -6048 -4519
rect -6041 -4522 -6017 -4518
rect -6010 -4522 -5991 -4518
rect -6121 -4528 -6059 -4526
rect -6114 -4530 -6059 -4528
rect -6041 -4533 -6037 -4522
rect -6010 -4525 -6006 -4522
rect -6018 -4539 -6014 -4535
rect -6024 -4540 -5999 -4539
rect -6024 -4544 -6004 -4540
rect -6024 -4545 -5999 -4544
rect -6060 -4557 -6056 -4553
rect -6060 -4561 -6044 -4557
rect -6057 -4601 -6034 -4597
rect -6053 -4603 -6034 -4601
rect -6057 -4612 -6053 -4607
rect -6038 -4612 -6034 -4603
rect -6021 -4608 -5997 -4607
rect -6021 -4612 -6005 -4608
rect -6001 -4612 -5997 -4608
rect -6021 -4614 -5997 -4612
rect -6015 -4619 -6011 -4614
rect -6046 -4640 -6042 -4632
rect -6046 -4644 -6034 -4640
rect -6038 -4646 -6034 -4644
rect -6007 -4646 -6003 -4639
rect -5979 -4646 -5972 -4511
rect -6130 -4651 -6045 -4647
rect -6038 -4650 -6014 -4646
rect -6007 -4650 -5972 -4646
rect -6136 -4655 -6056 -4654
rect -6136 -4658 -6134 -4655
rect -6128 -4658 -6056 -4655
rect -6038 -4661 -6034 -4650
rect -6007 -4653 -6003 -4650
rect -6015 -4667 -6011 -4663
rect -6021 -4668 -5996 -4667
rect -6021 -4672 -6001 -4668
rect -6021 -4673 -5996 -4672
rect -6057 -4685 -6053 -4681
rect -6057 -4689 -6041 -4685
rect -6055 -4721 -6032 -4717
rect -6051 -4723 -6032 -4721
rect -6055 -4732 -6051 -4727
rect -6036 -4732 -6032 -4723
rect -6019 -4728 -5995 -4727
rect -6019 -4732 -6003 -4728
rect -5999 -4732 -5995 -4728
rect -6019 -4734 -5995 -4732
rect -6013 -4739 -6009 -4734
rect -6044 -4760 -6040 -4752
rect -6044 -4764 -6032 -4760
rect -6036 -4766 -6032 -4764
rect -6005 -4766 -6001 -4759
rect -5956 -4766 -5951 -4610
rect -6122 -4771 -6043 -4767
rect -6036 -4770 -6012 -4766
rect -6005 -4770 -5951 -4766
rect -6128 -4776 -6054 -4774
rect -6122 -4778 -6054 -4776
rect -6036 -4781 -6032 -4770
rect -6005 -4773 -6001 -4770
rect -6013 -4787 -6009 -4783
rect -6019 -4788 -5994 -4787
rect -6019 -4792 -5999 -4788
rect -6019 -4793 -5994 -4792
rect -6055 -4805 -6051 -4801
rect -6055 -4809 -6039 -4805
rect -6053 -4862 -6030 -4858
rect -6049 -4864 -6030 -4862
rect -6053 -4873 -6049 -4868
rect -6034 -4873 -6030 -4864
rect -6017 -4869 -5993 -4868
rect -6017 -4873 -6001 -4869
rect -5997 -4873 -5993 -4869
rect -6017 -4875 -5993 -4873
rect -6011 -4880 -6007 -4875
rect -6042 -4901 -6038 -4893
rect -6042 -4905 -6030 -4901
rect -6034 -4907 -6030 -4905
rect -6003 -4907 -5999 -4900
rect -5937 -4907 -5932 -4669
rect -5078 -4717 -5074 -4269
rect -4914 -4291 -4910 -4269
rect -4906 -4717 -4902 -4391
rect -4740 -4324 -4736 -4269
rect -4732 -4717 -4728 -4424
rect -4616 -4395 -4612 -4269
rect -4608 -4717 -4604 -4495
rect -4477 -4494 -4473 -4050
rect -4398 -3956 -4393 -3365
rect -4286 -3398 -4282 -3389
rect -4286 -3403 -4285 -3398
rect -4286 -3407 -4282 -3403
rect -4294 -3437 -4290 -3427
rect -4293 -3470 -4289 -3467
rect -4299 -3474 -4298 -3470
rect -4294 -3474 -4289 -3470
rect -4293 -3480 -4289 -3474
rect -4285 -3530 -4281 -3520
rect -4285 -3535 -4284 -3530
rect -4285 -3538 -4281 -3535
rect -4293 -3568 -4289 -3558
rect -4293 -3601 -4289 -3598
rect -4299 -3605 -4298 -3601
rect -4294 -3605 -4289 -3601
rect -4293 -3611 -4289 -3605
rect -4285 -3660 -4281 -3651
rect -4285 -3665 -4284 -3660
rect -4285 -3669 -4281 -3665
rect -4293 -3699 -4289 -3689
rect -4294 -3744 -4290 -3741
rect -4300 -3748 -4299 -3744
rect -4295 -3748 -4290 -3744
rect -4294 -3754 -4290 -3748
rect -4286 -3803 -4282 -3794
rect -4286 -3808 -4285 -3803
rect -4286 -3812 -4282 -3808
rect -4294 -3842 -4290 -3832
rect -4209 -3853 -4204 -2947
rect -4148 -3710 -4143 -2902
rect -4046 -3582 -4041 -2813
rect -3944 -3452 -3939 -2752
rect -3891 -3278 -3886 -2658
rect -3734 -3187 -3706 -3184
rect -3733 -3193 -3730 -3187
rect -3709 -3188 -3706 -3187
rect -3709 -3191 -3638 -3188
rect -3756 -3215 -3747 -3214
rect -3752 -3217 -3747 -3215
rect -3742 -3216 -3732 -3213
rect -3724 -3213 -3721 -3205
rect -3694 -3197 -3691 -3191
rect -3675 -3197 -3672 -3191
rect -3724 -3216 -3703 -3213
rect -3724 -3219 -3721 -3216
rect -3733 -3229 -3730 -3225
rect -3739 -3231 -3715 -3229
rect -3739 -3232 -3721 -3231
rect -3716 -3232 -3715 -3231
rect -3706 -3239 -3703 -3216
rect -3665 -3197 -3645 -3194
rect -3665 -3203 -3662 -3197
rect -3648 -3203 -3645 -3197
rect -3684 -3224 -3681 -3221
rect -3684 -3227 -3666 -3224
rect -3526 -3218 -3514 -3214
rect -3400 -3215 -3390 -3211
rect -3310 -3218 -3298 -3214
rect -3184 -3215 -3174 -3211
rect -3656 -3234 -3653 -3227
rect -3564 -3229 -3539 -3225
rect -3479 -3229 -3454 -3225
rect -3412 -3226 -3387 -3222
rect -3558 -3233 -3554 -3229
rect -3473 -3233 -3469 -3229
rect -3412 -3230 -3408 -3226
rect -3391 -3230 -3387 -3226
rect -3656 -3237 -3639 -3234
rect -3734 -3240 -3715 -3239
rect -3739 -3242 -3715 -3240
rect -3706 -3242 -3663 -3239
rect -3733 -3248 -3730 -3242
rect -3642 -3249 -3639 -3237
rect -3550 -3249 -3546 -3241
rect -3515 -3249 -3511 -3241
rect -3677 -3253 -3652 -3250
rect -3642 -3253 -3557 -3249
rect -3550 -3253 -3511 -3249
rect -3677 -3255 -3674 -3253
rect -3784 -3271 -3747 -3268
rect -3742 -3271 -3732 -3268
rect -3724 -3268 -3721 -3260
rect -3712 -3258 -3674 -3255
rect -3642 -3256 -3639 -3253
rect -3712 -3268 -3709 -3258
rect -3671 -3259 -3639 -3256
rect -3671 -3262 -3668 -3259
rect -3724 -3271 -3709 -3268
rect -3724 -3274 -3721 -3271
rect -3891 -3284 -3806 -3278
rect -3672 -3265 -3666 -3262
rect -3733 -3284 -3730 -3280
rect -3712 -3281 -3707 -3278
rect -3694 -3278 -3691 -3274
rect -3647 -3278 -3644 -3274
rect -3702 -3281 -3638 -3278
rect -3712 -3284 -3709 -3281
rect -3739 -3287 -3709 -3284
rect -3633 -3292 -3629 -3253
rect -3550 -3256 -3546 -3253
rect -3515 -3257 -3511 -3253
rect -3558 -3264 -3554 -3260
rect -3383 -3226 -3370 -3222
rect -3383 -3230 -3379 -3226
rect -3348 -3229 -3323 -3225
rect -3263 -3229 -3238 -3225
rect -3196 -3226 -3171 -3222
rect -3342 -3233 -3338 -3229
rect -3257 -3233 -3253 -3229
rect -3196 -3230 -3192 -3226
rect -3175 -3230 -3171 -3226
rect -3507 -3249 -3503 -3241
rect -3465 -3249 -3461 -3241
rect -3404 -3249 -3400 -3238
rect -3334 -3249 -3330 -3241
rect -3299 -3249 -3295 -3241
rect -3507 -3253 -3472 -3249
rect -3465 -3253 -3411 -3249
rect -3404 -3253 -3341 -3249
rect -3334 -3253 -3295 -3249
rect -3507 -3257 -3503 -3253
rect -3465 -3256 -3461 -3253
rect -3404 -3259 -3400 -3253
rect -3334 -3256 -3330 -3253
rect -3473 -3264 -3469 -3260
rect -3564 -3267 -3539 -3264
rect -3479 -3267 -3454 -3264
rect -3412 -3268 -3408 -3263
rect -3391 -3268 -3387 -3263
rect -3528 -3275 -3514 -3271
rect -3412 -3272 -3387 -3268
rect -3383 -3268 -3379 -3263
rect -3299 -3257 -3295 -3253
rect -3342 -3264 -3338 -3260
rect -3167 -3226 -3154 -3222
rect -3167 -3230 -3163 -3226
rect -3291 -3249 -3287 -3241
rect -3249 -3249 -3245 -3241
rect -3188 -3249 -3184 -3238
rect -3291 -3253 -3256 -3249
rect -3249 -3253 -3195 -3249
rect -3188 -3253 -3148 -3249
rect -3291 -3257 -3287 -3253
rect -3249 -3256 -3245 -3253
rect -3188 -3259 -3184 -3253
rect -3257 -3264 -3253 -3260
rect -3348 -3267 -3323 -3264
rect -3263 -3267 -3238 -3264
rect -3196 -3268 -3192 -3263
rect -3175 -3268 -3171 -3263
rect -3383 -3272 -3370 -3268
rect -3312 -3275 -3298 -3271
rect -3196 -3272 -3171 -3268
rect -3167 -3268 -3163 -3263
rect -3167 -3272 -3154 -3268
rect -3528 -3278 -3524 -3275
rect -3399 -3279 -3390 -3275
rect -3183 -3279 -3174 -3275
rect -3803 -3371 -3775 -3368
rect -3802 -3377 -3799 -3371
rect -3778 -3372 -3775 -3371
rect -3778 -3375 -3707 -3372
rect -3829 -3401 -3816 -3398
rect -3811 -3400 -3801 -3397
rect -3793 -3397 -3790 -3389
rect -3763 -3381 -3760 -3375
rect -3744 -3381 -3741 -3375
rect -3793 -3400 -3772 -3397
rect -3793 -3403 -3790 -3400
rect -3802 -3413 -3799 -3409
rect -3808 -3415 -3784 -3413
rect -3808 -3416 -3790 -3415
rect -3785 -3416 -3784 -3415
rect -3775 -3423 -3772 -3400
rect -3734 -3381 -3714 -3378
rect -3734 -3387 -3731 -3381
rect -3717 -3387 -3714 -3381
rect -3753 -3408 -3750 -3405
rect -3753 -3411 -3735 -3408
rect -3531 -3402 -3519 -3398
rect -3405 -3399 -3395 -3395
rect -3315 -3402 -3303 -3398
rect -3189 -3399 -3179 -3395
rect -3725 -3418 -3722 -3411
rect -3569 -3413 -3544 -3409
rect -3484 -3413 -3459 -3409
rect -3417 -3410 -3392 -3406
rect -3563 -3417 -3559 -3413
rect -3478 -3417 -3474 -3413
rect -3417 -3414 -3413 -3410
rect -3396 -3414 -3392 -3410
rect -3725 -3421 -3708 -3418
rect -3803 -3424 -3784 -3423
rect -3808 -3426 -3784 -3424
rect -3775 -3426 -3732 -3423
rect -3802 -3432 -3799 -3426
rect -3711 -3432 -3708 -3421
rect -3711 -3433 -3698 -3432
rect -3555 -3433 -3551 -3425
rect -3520 -3433 -3516 -3425
rect -3746 -3437 -3721 -3434
rect -3711 -3436 -3562 -3433
rect -3746 -3439 -3743 -3437
rect -3944 -3455 -3816 -3452
rect -3811 -3455 -3801 -3452
rect -3793 -3452 -3790 -3444
rect -3781 -3442 -3743 -3439
rect -3711 -3440 -3708 -3436
rect -3781 -3452 -3778 -3442
rect -3740 -3443 -3708 -3440
rect -3702 -3437 -3562 -3436
rect -3555 -3437 -3516 -3433
rect -3740 -3446 -3737 -3443
rect -3793 -3455 -3778 -3452
rect -3793 -3458 -3790 -3455
rect -3741 -3449 -3735 -3446
rect -3802 -3468 -3799 -3464
rect -3781 -3465 -3776 -3462
rect -3763 -3462 -3760 -3458
rect -3716 -3462 -3713 -3458
rect -3771 -3465 -3707 -3462
rect -3781 -3468 -3778 -3465
rect -3808 -3471 -3778 -3468
rect -3702 -3476 -3698 -3437
rect -3555 -3440 -3551 -3437
rect -3520 -3441 -3516 -3437
rect -3563 -3448 -3559 -3444
rect -3388 -3410 -3375 -3406
rect -3388 -3414 -3384 -3410
rect -3353 -3413 -3328 -3409
rect -3268 -3413 -3243 -3409
rect -3201 -3410 -3176 -3406
rect -3347 -3417 -3343 -3413
rect -3262 -3417 -3258 -3413
rect -3201 -3414 -3197 -3410
rect -3180 -3414 -3176 -3410
rect -3512 -3433 -3508 -3425
rect -3470 -3433 -3466 -3425
rect -3409 -3433 -3405 -3422
rect -3339 -3433 -3335 -3425
rect -3304 -3433 -3300 -3425
rect -3512 -3437 -3477 -3433
rect -3470 -3437 -3416 -3433
rect -3409 -3437 -3346 -3433
rect -3339 -3437 -3300 -3433
rect -3512 -3441 -3508 -3437
rect -3470 -3440 -3466 -3437
rect -3409 -3443 -3405 -3437
rect -3339 -3440 -3335 -3437
rect -3478 -3448 -3474 -3444
rect -3569 -3451 -3544 -3448
rect -3484 -3451 -3459 -3448
rect -3417 -3452 -3413 -3447
rect -3396 -3452 -3392 -3447
rect -3533 -3459 -3519 -3455
rect -3417 -3456 -3392 -3452
rect -3388 -3452 -3384 -3447
rect -3304 -3441 -3300 -3437
rect -3347 -3448 -3343 -3444
rect -3172 -3410 -3159 -3406
rect -3172 -3414 -3168 -3410
rect -3296 -3433 -3292 -3425
rect -3254 -3433 -3250 -3425
rect -3193 -3433 -3189 -3422
rect -3296 -3437 -3261 -3433
rect -3254 -3437 -3200 -3433
rect -3193 -3437 -3153 -3433
rect -3296 -3441 -3292 -3437
rect -3254 -3440 -3250 -3437
rect -3193 -3443 -3189 -3437
rect -3262 -3448 -3258 -3444
rect -3353 -3451 -3328 -3448
rect -3268 -3451 -3243 -3448
rect -3201 -3452 -3197 -3447
rect -3180 -3452 -3176 -3447
rect -3388 -3456 -3375 -3452
rect -3317 -3459 -3303 -3455
rect -3201 -3456 -3176 -3452
rect -3172 -3452 -3168 -3447
rect -3172 -3456 -3159 -3452
rect -3533 -3462 -3529 -3459
rect -3404 -3463 -3395 -3459
rect -3188 -3463 -3179 -3459
rect -3808 -3501 -3780 -3498
rect -3807 -3507 -3804 -3501
rect -3783 -3502 -3780 -3501
rect -3783 -3505 -3712 -3502
rect -3831 -3530 -3821 -3528
rect -3826 -3531 -3821 -3530
rect -3816 -3530 -3806 -3527
rect -3798 -3527 -3795 -3519
rect -3768 -3511 -3765 -3505
rect -3749 -3511 -3746 -3505
rect -3798 -3530 -3777 -3527
rect -3798 -3533 -3795 -3530
rect -3807 -3543 -3804 -3539
rect -3813 -3545 -3789 -3543
rect -3813 -3546 -3795 -3545
rect -3790 -3546 -3789 -3545
rect -3780 -3553 -3777 -3530
rect -3739 -3511 -3719 -3508
rect -3739 -3517 -3736 -3511
rect -3722 -3517 -3719 -3511
rect -3758 -3538 -3755 -3535
rect -3758 -3541 -3740 -3538
rect -3534 -3533 -3522 -3529
rect -3408 -3530 -3398 -3526
rect -3318 -3533 -3306 -3529
rect -3192 -3530 -3182 -3526
rect -3730 -3548 -3727 -3541
rect -3572 -3544 -3547 -3540
rect -3487 -3544 -3462 -3540
rect -3420 -3541 -3395 -3537
rect -3566 -3548 -3562 -3544
rect -3481 -3548 -3477 -3544
rect -3420 -3545 -3416 -3541
rect -3399 -3545 -3395 -3541
rect -3730 -3551 -3713 -3548
rect -3808 -3554 -3789 -3553
rect -3813 -3556 -3789 -3554
rect -3780 -3556 -3737 -3553
rect -3807 -3562 -3804 -3556
rect -3716 -3562 -3713 -3551
rect -3751 -3567 -3726 -3564
rect -3716 -3564 -3703 -3562
rect -3558 -3564 -3554 -3556
rect -3523 -3564 -3519 -3556
rect -3716 -3566 -3565 -3564
rect -3751 -3569 -3748 -3567
rect -4046 -3585 -3821 -3582
rect -3816 -3585 -3806 -3582
rect -3798 -3582 -3795 -3574
rect -3786 -3572 -3748 -3569
rect -3716 -3570 -3713 -3566
rect -3786 -3582 -3783 -3572
rect -3745 -3573 -3713 -3570
rect -3707 -3568 -3565 -3566
rect -3558 -3568 -3519 -3564
rect -3745 -3576 -3742 -3573
rect -3798 -3585 -3783 -3582
rect -3798 -3588 -3795 -3585
rect -3746 -3579 -3740 -3576
rect -3807 -3598 -3804 -3594
rect -3786 -3595 -3781 -3592
rect -3768 -3592 -3765 -3588
rect -3721 -3592 -3718 -3588
rect -3776 -3595 -3712 -3592
rect -3786 -3598 -3783 -3595
rect -3813 -3601 -3783 -3598
rect -3707 -3606 -3703 -3568
rect -3558 -3571 -3554 -3568
rect -3523 -3572 -3519 -3568
rect -3566 -3579 -3562 -3575
rect -3391 -3541 -3378 -3537
rect -3391 -3545 -3387 -3541
rect -3356 -3544 -3331 -3540
rect -3271 -3544 -3246 -3540
rect -3204 -3541 -3179 -3537
rect -3350 -3548 -3346 -3544
rect -3265 -3548 -3261 -3544
rect -3204 -3545 -3200 -3541
rect -3183 -3545 -3179 -3541
rect -3515 -3564 -3511 -3556
rect -3473 -3564 -3469 -3556
rect -3412 -3564 -3408 -3553
rect -3342 -3564 -3338 -3556
rect -3307 -3564 -3303 -3556
rect -3515 -3568 -3480 -3564
rect -3473 -3568 -3419 -3564
rect -3412 -3568 -3349 -3564
rect -3342 -3568 -3303 -3564
rect -3515 -3572 -3511 -3568
rect -3473 -3571 -3469 -3568
rect -3412 -3574 -3408 -3568
rect -3342 -3571 -3338 -3568
rect -3481 -3579 -3477 -3575
rect -3572 -3582 -3547 -3579
rect -3487 -3582 -3462 -3579
rect -3420 -3583 -3416 -3578
rect -3399 -3583 -3395 -3578
rect -3536 -3590 -3522 -3586
rect -3420 -3587 -3395 -3583
rect -3391 -3583 -3387 -3578
rect -3307 -3572 -3303 -3568
rect -3350 -3579 -3346 -3575
rect -3175 -3541 -3162 -3537
rect -3175 -3545 -3171 -3541
rect -3299 -3564 -3295 -3556
rect -3257 -3564 -3253 -3556
rect -3196 -3564 -3192 -3553
rect -3299 -3568 -3264 -3564
rect -3257 -3568 -3203 -3564
rect -3196 -3568 -3156 -3564
rect -3299 -3572 -3295 -3568
rect -3257 -3571 -3253 -3568
rect -3196 -3574 -3192 -3568
rect -3265 -3579 -3261 -3575
rect -3356 -3582 -3331 -3579
rect -3271 -3582 -3246 -3579
rect -3204 -3583 -3200 -3578
rect -3183 -3583 -3179 -3578
rect -3391 -3587 -3378 -3583
rect -3320 -3590 -3306 -3586
rect -3204 -3587 -3179 -3583
rect -3175 -3583 -3171 -3578
rect -3175 -3587 -3162 -3583
rect -3536 -3593 -3532 -3590
rect -3407 -3594 -3398 -3590
rect -3191 -3594 -3182 -3590
rect -3804 -3629 -3776 -3626
rect -3803 -3635 -3800 -3629
rect -3779 -3630 -3776 -3629
rect -3779 -3633 -3708 -3630
rect -3829 -3659 -3817 -3656
rect -3829 -3660 -3824 -3659
rect -3812 -3658 -3802 -3655
rect -3794 -3655 -3791 -3647
rect -3764 -3639 -3761 -3633
rect -3745 -3639 -3742 -3633
rect -3794 -3658 -3773 -3655
rect -3794 -3661 -3791 -3658
rect -3803 -3671 -3800 -3667
rect -3809 -3673 -3785 -3671
rect -3809 -3674 -3791 -3673
rect -3786 -3674 -3785 -3673
rect -3776 -3681 -3773 -3658
rect -3735 -3639 -3715 -3636
rect -3735 -3645 -3732 -3639
rect -3718 -3645 -3715 -3639
rect -3754 -3666 -3751 -3663
rect -3754 -3669 -3736 -3666
rect -3547 -3663 -3535 -3659
rect -3421 -3660 -3411 -3656
rect -3331 -3663 -3319 -3659
rect -3205 -3660 -3195 -3656
rect -3726 -3676 -3723 -3669
rect -3585 -3674 -3560 -3670
rect -3500 -3674 -3475 -3670
rect -3433 -3671 -3408 -3667
rect -3726 -3679 -3709 -3676
rect -3804 -3682 -3785 -3681
rect -3809 -3684 -3785 -3682
rect -3776 -3684 -3733 -3681
rect -3803 -3690 -3800 -3684
rect -3712 -3690 -3709 -3679
rect -3579 -3678 -3575 -3674
rect -3494 -3678 -3490 -3674
rect -3433 -3675 -3429 -3671
rect -3412 -3675 -3408 -3671
rect -3747 -3695 -3722 -3692
rect -3712 -3694 -3699 -3690
rect -3571 -3694 -3567 -3686
rect -3536 -3694 -3532 -3686
rect -3747 -3697 -3744 -3695
rect -4148 -3713 -3817 -3710
rect -3812 -3713 -3802 -3710
rect -3794 -3710 -3791 -3702
rect -3782 -3700 -3744 -3697
rect -3712 -3698 -3709 -3694
rect -3782 -3710 -3779 -3700
rect -3741 -3701 -3709 -3698
rect -3703 -3698 -3578 -3694
rect -3571 -3698 -3532 -3694
rect -3741 -3704 -3738 -3701
rect -3794 -3713 -3779 -3710
rect -3794 -3716 -3791 -3713
rect -3742 -3707 -3736 -3704
rect -3803 -3726 -3800 -3722
rect -3782 -3723 -3777 -3720
rect -3764 -3720 -3761 -3716
rect -3717 -3720 -3714 -3716
rect -3772 -3723 -3708 -3720
rect -3782 -3726 -3779 -3723
rect -3809 -3729 -3779 -3726
rect -3703 -3734 -3699 -3698
rect -3571 -3701 -3567 -3698
rect -3536 -3702 -3532 -3698
rect -3579 -3709 -3575 -3705
rect -3404 -3671 -3391 -3667
rect -3404 -3675 -3400 -3671
rect -3369 -3674 -3344 -3670
rect -3284 -3674 -3259 -3670
rect -3217 -3671 -3192 -3667
rect -3363 -3678 -3359 -3674
rect -3278 -3678 -3274 -3674
rect -3217 -3675 -3213 -3671
rect -3196 -3675 -3192 -3671
rect -3528 -3694 -3524 -3686
rect -3486 -3694 -3482 -3686
rect -3425 -3694 -3421 -3683
rect -3355 -3694 -3351 -3686
rect -3320 -3694 -3316 -3686
rect -3528 -3698 -3493 -3694
rect -3486 -3698 -3432 -3694
rect -3425 -3698 -3362 -3694
rect -3355 -3698 -3316 -3694
rect -3528 -3702 -3524 -3698
rect -3486 -3701 -3482 -3698
rect -3425 -3704 -3421 -3698
rect -3355 -3701 -3351 -3698
rect -3494 -3709 -3490 -3705
rect -3585 -3712 -3560 -3709
rect -3500 -3712 -3475 -3709
rect -3433 -3713 -3429 -3708
rect -3412 -3713 -3408 -3708
rect -3549 -3720 -3535 -3716
rect -3433 -3717 -3408 -3713
rect -3404 -3713 -3400 -3708
rect -3320 -3702 -3316 -3698
rect -3363 -3709 -3359 -3705
rect -3188 -3671 -3175 -3667
rect -3188 -3675 -3184 -3671
rect -3312 -3694 -3308 -3686
rect -3270 -3694 -3266 -3686
rect -3209 -3694 -3205 -3683
rect -3312 -3698 -3277 -3694
rect -3270 -3698 -3216 -3694
rect -3209 -3698 -3169 -3694
rect -3312 -3702 -3308 -3698
rect -3270 -3701 -3266 -3698
rect -3209 -3704 -3205 -3698
rect -3278 -3709 -3274 -3705
rect -3369 -3712 -3344 -3709
rect -3284 -3712 -3259 -3709
rect -3217 -3713 -3213 -3708
rect -3196 -3713 -3192 -3708
rect -3404 -3717 -3391 -3713
rect -3333 -3720 -3319 -3716
rect -3217 -3717 -3192 -3713
rect -3188 -3713 -3184 -3708
rect -3188 -3717 -3175 -3713
rect -3549 -3723 -3545 -3720
rect -3420 -3724 -3411 -3720
rect -3204 -3724 -3195 -3720
rect -3803 -3772 -3775 -3769
rect -3802 -3778 -3799 -3772
rect -3778 -3773 -3775 -3772
rect -3778 -3776 -3707 -3773
rect -3828 -3802 -3816 -3799
rect -3828 -3803 -3823 -3802
rect -3811 -3801 -3801 -3798
rect -3793 -3798 -3790 -3790
rect -3763 -3782 -3760 -3776
rect -3744 -3782 -3741 -3776
rect -3793 -3801 -3772 -3798
rect -3793 -3804 -3790 -3801
rect -3802 -3814 -3799 -3810
rect -3808 -3816 -3784 -3814
rect -3808 -3817 -3790 -3816
rect -3785 -3817 -3784 -3816
rect -3775 -3824 -3772 -3801
rect -3734 -3782 -3714 -3779
rect -3734 -3788 -3731 -3782
rect -3717 -3788 -3714 -3782
rect -3753 -3809 -3750 -3806
rect -3753 -3812 -3735 -3809
rect -3546 -3806 -3534 -3802
rect -3420 -3803 -3410 -3799
rect -3330 -3806 -3318 -3802
rect -3204 -3803 -3194 -3799
rect -3725 -3819 -3722 -3812
rect -3584 -3817 -3559 -3813
rect -3499 -3817 -3474 -3813
rect -3432 -3814 -3407 -3810
rect -3725 -3822 -3708 -3819
rect -3803 -3825 -3784 -3824
rect -3808 -3827 -3784 -3825
rect -3775 -3827 -3732 -3824
rect -3802 -3833 -3799 -3827
rect -3711 -3833 -3708 -3822
rect -3578 -3821 -3574 -3817
rect -3493 -3821 -3489 -3817
rect -3432 -3818 -3428 -3814
rect -3411 -3818 -3407 -3814
rect -3746 -3838 -3721 -3835
rect -3711 -3837 -3698 -3833
rect -3570 -3837 -3566 -3829
rect -3535 -3837 -3531 -3829
rect -3746 -3840 -3743 -3838
rect -4209 -3856 -3816 -3853
rect -3811 -3856 -3801 -3853
rect -3793 -3853 -3790 -3845
rect -3781 -3843 -3743 -3840
rect -3711 -3841 -3708 -3837
rect -3781 -3853 -3778 -3843
rect -3740 -3844 -3708 -3841
rect -3702 -3841 -3577 -3837
rect -3570 -3841 -3531 -3837
rect -3740 -3847 -3737 -3844
rect -3793 -3856 -3778 -3853
rect -3793 -3859 -3790 -3856
rect -3741 -3850 -3735 -3847
rect -3802 -3869 -3799 -3865
rect -3781 -3866 -3776 -3863
rect -3763 -3863 -3760 -3859
rect -3716 -3863 -3713 -3859
rect -3771 -3866 -3707 -3863
rect -3781 -3869 -3778 -3866
rect -3808 -3872 -3778 -3869
rect -3702 -3877 -3698 -3841
rect -3570 -3844 -3566 -3841
rect -3535 -3845 -3531 -3841
rect -3578 -3852 -3574 -3848
rect -3403 -3814 -3390 -3810
rect -3403 -3818 -3399 -3814
rect -3368 -3817 -3343 -3813
rect -3283 -3817 -3258 -3813
rect -3216 -3814 -3191 -3810
rect -3362 -3821 -3358 -3817
rect -3277 -3821 -3273 -3817
rect -3216 -3818 -3212 -3814
rect -3195 -3818 -3191 -3814
rect -3527 -3837 -3523 -3829
rect -3485 -3837 -3481 -3829
rect -3424 -3837 -3420 -3826
rect -3354 -3837 -3350 -3829
rect -3319 -3837 -3315 -3829
rect -3527 -3841 -3492 -3837
rect -3485 -3841 -3431 -3837
rect -3424 -3841 -3361 -3837
rect -3354 -3841 -3315 -3837
rect -3527 -3845 -3523 -3841
rect -3485 -3844 -3481 -3841
rect -3424 -3847 -3420 -3841
rect -3354 -3844 -3350 -3841
rect -3493 -3852 -3489 -3848
rect -3584 -3855 -3559 -3852
rect -3499 -3855 -3474 -3852
rect -3432 -3856 -3428 -3851
rect -3411 -3856 -3407 -3851
rect -3548 -3863 -3534 -3859
rect -3432 -3860 -3407 -3856
rect -3403 -3856 -3399 -3851
rect -3319 -3845 -3315 -3841
rect -3362 -3852 -3358 -3848
rect -3187 -3814 -3174 -3810
rect -3187 -3818 -3183 -3814
rect -3311 -3837 -3307 -3829
rect -3269 -3837 -3265 -3829
rect -3208 -3837 -3204 -3826
rect -3311 -3841 -3276 -3837
rect -3269 -3841 -3215 -3837
rect -3208 -3841 -3168 -3837
rect -3311 -3845 -3307 -3841
rect -3269 -3844 -3265 -3841
rect -3208 -3847 -3204 -3841
rect -3277 -3852 -3273 -3848
rect -3368 -3855 -3343 -3852
rect -3283 -3855 -3258 -3852
rect -3216 -3856 -3212 -3851
rect -3195 -3856 -3191 -3851
rect -3403 -3860 -3390 -3856
rect -3332 -3863 -3318 -3859
rect -3216 -3860 -3191 -3856
rect -3187 -3856 -3183 -3851
rect -3187 -3860 -3174 -3856
rect -3548 -3866 -3544 -3863
rect -3419 -3867 -3410 -3863
rect -3203 -3867 -3194 -3863
rect -4294 -3896 -4290 -3893
rect -4300 -3900 -4299 -3896
rect -4295 -3900 -4290 -3896
rect -4294 -3906 -4290 -3900
rect -3561 -3924 -3549 -3920
rect -3435 -3921 -3425 -3917
rect -3345 -3924 -3333 -3920
rect -3219 -3921 -3209 -3917
rect -3599 -3935 -3574 -3931
rect -3514 -3935 -3489 -3931
rect -3447 -3932 -3422 -3928
rect -4286 -3955 -4282 -3946
rect -3593 -3939 -3589 -3935
rect -3508 -3939 -3504 -3935
rect -3447 -3936 -3443 -3932
rect -3426 -3936 -3422 -3932
rect -3585 -3955 -3581 -3947
rect -3550 -3955 -3546 -3947
rect -4286 -3960 -4285 -3955
rect -3605 -3959 -3592 -3955
rect -3585 -3959 -3546 -3955
rect -4469 -4717 -4465 -4594
rect -4398 -4553 -4394 -3961
rect -4286 -3964 -4282 -3960
rect -3585 -3962 -3581 -3959
rect -3550 -3963 -3546 -3959
rect -3593 -3970 -3589 -3966
rect -3418 -3932 -3405 -3928
rect -3418 -3936 -3414 -3932
rect -3383 -3935 -3358 -3931
rect -3298 -3935 -3273 -3931
rect -3231 -3932 -3206 -3928
rect -3377 -3939 -3373 -3935
rect -3292 -3939 -3288 -3935
rect -3231 -3936 -3227 -3932
rect -3210 -3936 -3206 -3932
rect -3542 -3955 -3538 -3947
rect -3500 -3955 -3496 -3947
rect -3439 -3955 -3435 -3944
rect -3369 -3955 -3365 -3947
rect -3334 -3955 -3330 -3947
rect -3542 -3959 -3507 -3955
rect -3500 -3959 -3446 -3955
rect -3439 -3959 -3376 -3955
rect -3369 -3959 -3330 -3955
rect -3542 -3963 -3538 -3959
rect -3500 -3962 -3496 -3959
rect -3439 -3965 -3435 -3959
rect -3369 -3962 -3365 -3959
rect -3508 -3970 -3504 -3966
rect -3599 -3973 -3574 -3970
rect -3514 -3973 -3489 -3970
rect -3447 -3974 -3443 -3969
rect -3426 -3974 -3422 -3969
rect -3563 -3981 -3549 -3977
rect -3447 -3978 -3422 -3974
rect -3418 -3974 -3414 -3969
rect -3334 -3963 -3330 -3959
rect -3377 -3970 -3373 -3966
rect -3202 -3932 -3189 -3928
rect -3202 -3936 -3198 -3932
rect -3326 -3955 -3322 -3947
rect -3284 -3955 -3280 -3947
rect -3223 -3955 -3219 -3944
rect -3326 -3959 -3291 -3955
rect -3284 -3959 -3230 -3955
rect -3223 -3959 -3183 -3955
rect -3326 -3963 -3322 -3959
rect -3284 -3962 -3280 -3959
rect -3223 -3965 -3219 -3959
rect -3292 -3970 -3288 -3966
rect -3383 -3973 -3358 -3970
rect -3298 -3973 -3273 -3970
rect -3231 -3974 -3227 -3969
rect -3210 -3974 -3206 -3969
rect -3418 -3978 -3405 -3974
rect -3347 -3981 -3333 -3977
rect -3231 -3978 -3206 -3974
rect -3202 -3974 -3198 -3969
rect -3202 -3978 -3189 -3974
rect -3563 -3984 -3559 -3981
rect -4294 -3994 -4290 -3984
rect -3434 -3985 -3425 -3981
rect -3218 -3985 -3209 -3981
rect -5078 -4718 -4465 -4717
rect -4390 -4718 -4386 -4653
rect -5078 -4722 -4386 -4718
rect -5078 -4811 -5074 -4722
rect -5231 -4862 -5227 -4859
rect -5237 -4866 -5236 -4862
rect -5232 -4866 -5227 -4862
rect -6120 -4912 -6041 -4908
rect -6034 -4911 -6010 -4907
rect -6003 -4911 -5932 -4907
rect -5231 -4872 -5227 -4866
rect -6126 -4917 -6052 -4915
rect -6120 -4919 -6052 -4917
rect -6034 -4922 -6030 -4911
rect -6003 -4914 -5999 -4911
rect -5223 -4922 -5219 -4912
rect -5070 -4920 -5066 -4911
rect -6011 -4928 -6007 -4924
rect -5223 -4927 -5086 -4922
rect -6017 -4929 -5992 -4928
rect -6017 -4933 -5997 -4929
rect -5223 -4930 -5219 -4927
rect -6017 -4934 -5992 -4933
rect -6053 -4946 -6049 -4942
rect -6053 -4950 -6037 -4946
rect -5231 -4960 -5227 -4950
<< m2contact >>
rect -5882 -2602 -5877 -2595
rect -8122 -3048 -8117 -3043
rect -7704 -3041 -7699 -3036
rect -7980 -3054 -7975 -3049
rect -7838 -3052 -7833 -3047
rect -7569 -3051 -7564 -3046
rect -6091 -3477 -6086 -3472
rect -6276 -3532 -6271 -3527
rect -6091 -3531 -6086 -3526
rect -5977 -3515 -5972 -3510
rect -5984 -3604 -5979 -3599
rect -6098 -3649 -6093 -3644
rect -6185 -3704 -6180 -3699
rect -6098 -3703 -6093 -3698
rect -6095 -3793 -6090 -3788
rect -5765 -2666 -5760 -2659
rect -5765 -3515 -5760 -3510
rect -5708 -2752 -5703 -2745
rect -3944 -2752 -3939 -2746
rect -5708 -3604 -5703 -3599
rect -5616 -2813 -5611 -2806
rect -5882 -3783 -5877 -3778
rect -6183 -3848 -6178 -3843
rect -6095 -3847 -6090 -3842
rect -5981 -3838 -5976 -3833
rect -4046 -2813 -4041 -2807
rect -5616 -3838 -5611 -3833
rect -5487 -2902 -5482 -2895
rect -4148 -2902 -4143 -2895
rect -5985 -3869 -5980 -3864
rect -5487 -3869 -5482 -3864
rect -5327 -2947 -5322 -2942
rect -6099 -3941 -6094 -3936
rect -6179 -3996 -6174 -3991
rect -6099 -3995 -6094 -3990
rect -4209 -2947 -4204 -2942
rect -5115 -3290 -5108 -3284
rect -4942 -3291 -4937 -3285
rect -4997 -3404 -4992 -3399
rect -4768 -3291 -4762 -3285
rect -4644 -3292 -4639 -3286
rect -5960 -4032 -5955 -4027
rect -5327 -4032 -5322 -4027
rect -6074 -4157 -6069 -4152
rect -6154 -4212 -6149 -4207
rect -6074 -4211 -6069 -4206
rect -4814 -3535 -4809 -3530
rect -4657 -3666 -4652 -3661
rect -4504 -3295 -4499 -3289
rect -4540 -3809 -4535 -3804
rect -5990 -4407 -5984 -4402
rect -6213 -4414 -6208 -4409
rect -6219 -4423 -6213 -4418
rect -5996 -4440 -5991 -4435
rect -6121 -4523 -6115 -4518
rect -5979 -4511 -5972 -4506
rect -6121 -4534 -6114 -4528
rect -6136 -4651 -6130 -4646
rect -5956 -4610 -5951 -4605
rect -6134 -4660 -6128 -4655
rect -6128 -4771 -6122 -4765
rect -5937 -4669 -5932 -4664
rect -6128 -4781 -6122 -4776
rect -6126 -4912 -6120 -4906
rect -4285 -3403 -4280 -3398
rect -4284 -3535 -4279 -3530
rect -4284 -3665 -4279 -3660
rect -4285 -3808 -4280 -3803
rect -3758 -3220 -3752 -3215
rect -3747 -3218 -3742 -3213
rect -3789 -3273 -3784 -3268
rect -3747 -3272 -3742 -3267
rect -3806 -3284 -3799 -3278
rect -3834 -3403 -3829 -3398
rect -3816 -3402 -3811 -3397
rect -3816 -3456 -3811 -3451
rect -3831 -3535 -3826 -3530
rect -3821 -3532 -3816 -3527
rect -3821 -3586 -3816 -3581
rect -3817 -3660 -3812 -3655
rect -3829 -3665 -3824 -3660
rect -3817 -3714 -3812 -3709
rect -3816 -3803 -3811 -3798
rect -3828 -3808 -3823 -3803
rect -3816 -3857 -3811 -3852
rect -4398 -3961 -4393 -3956
rect -4285 -3960 -4280 -3955
rect -3610 -3960 -3605 -3955
rect -6126 -4922 -6120 -4917
rect -5086 -4927 -5081 -4922
<< pm12contact >>
rect -6035 -3494 -6030 -3489
rect -6026 -3495 -6021 -3490
rect -6042 -3666 -6037 -3661
rect -6033 -3667 -6028 -3662
rect -6039 -3810 -6034 -3805
rect -6030 -3811 -6025 -3806
rect -6043 -3958 -6038 -3953
rect -6034 -3959 -6029 -3954
rect -5237 -3045 -5232 -3040
rect -5104 -3290 -5098 -3284
rect -4932 -3291 -4926 -3285
rect -5095 -3515 -5090 -3510
rect -4758 -3291 -4752 -3285
rect -4634 -3292 -4628 -3286
rect -4923 -3604 -4918 -3599
rect -5087 -3783 -5082 -3778
rect -6018 -4174 -6013 -4169
rect -6009 -4175 -6004 -4170
rect -4749 -3838 -4744 -3833
rect -4494 -3295 -4488 -3289
rect -4625 -3869 -4620 -3864
rect -4485 -4032 -4480 -4027
rect -4914 -4407 -4909 -4402
rect -4740 -4440 -4735 -4435
rect -4616 -4511 -4611 -4506
rect -4294 -3404 -4289 -3399
rect -4293 -3535 -4288 -3530
rect -4293 -3666 -4288 -3661
rect -4294 -3809 -4289 -3804
rect -3691 -3235 -3686 -3230
rect -3682 -3236 -3677 -3231
rect -3760 -3419 -3755 -3414
rect -3751 -3420 -3746 -3415
rect -3765 -3549 -3760 -3544
rect -3756 -3550 -3751 -3545
rect -3761 -3677 -3756 -3672
rect -3752 -3678 -3747 -3673
rect -3760 -3820 -3755 -3815
rect -3751 -3821 -3746 -3816
rect -4294 -3961 -4289 -3956
rect -4477 -4610 -4472 -4605
rect -4398 -4669 -4393 -4664
rect -5231 -4927 -5226 -4922
rect -5078 -4927 -5073 -4922
<< metal2 >>
rect -5877 -2596 -4685 -2595
rect -5877 -2602 -3839 -2596
rect -5760 -2660 -4304 -2659
rect -5760 -2666 -3887 -2660
rect -5703 -2746 -4319 -2745
rect -5703 -2752 -3944 -2746
rect -5611 -2807 -4242 -2806
rect -5611 -2813 -4046 -2807
rect -5482 -2902 -4148 -2895
rect -5322 -2947 -4209 -2942
rect -8122 -4207 -8118 -3048
rect -7980 -3049 -7976 -3042
rect -7980 -3991 -7976 -3054
rect -7838 -3843 -7833 -3052
rect -7704 -3699 -7699 -3041
rect -7569 -3046 -7565 -3039
rect -5240 -3045 -5237 -3040
rect -7569 -3527 -7565 -3051
rect -3844 -3214 -3839 -2602
rect -3844 -3215 -3756 -3214
rect -3844 -3220 -3758 -3215
rect -3746 -3224 -3743 -3218
rect -3746 -3227 -3709 -3224
rect -3712 -3230 -3709 -3227
rect -3712 -3233 -3691 -3230
rect -3682 -3246 -3679 -3236
rect -3745 -3249 -3679 -3246
rect -3745 -3267 -3742 -3249
rect -3789 -3278 -3784 -3273
rect -3799 -3284 -3784 -3278
rect -5108 -3290 -5104 -3284
rect -4937 -3291 -4932 -3285
rect -4762 -3291 -4758 -3285
rect -4639 -3292 -4634 -3286
rect -4499 -3295 -4494 -3289
rect -4992 -3404 -4294 -3399
rect -4280 -3403 -3834 -3398
rect -3815 -3408 -3812 -3402
rect -3815 -3411 -3778 -3408
rect -3781 -3414 -3778 -3411
rect -3781 -3417 -3760 -3414
rect -3751 -3430 -3748 -3420
rect -3814 -3433 -3748 -3430
rect -3814 -3451 -3811 -3433
rect -6090 -3483 -6087 -3477
rect -6090 -3486 -6053 -3483
rect -6056 -3489 -6053 -3486
rect -6056 -3492 -6035 -3489
rect -6026 -3505 -6023 -3495
rect -6089 -3508 -6023 -3505
rect -6089 -3526 -6086 -3508
rect -5972 -3515 -5765 -3510
rect -5760 -3515 -5095 -3510
rect -7569 -3532 -6388 -3527
rect -6383 -3532 -6276 -3527
rect -4809 -3535 -4293 -3530
rect -4279 -3535 -3831 -3530
rect -3820 -3538 -3817 -3532
rect -3820 -3541 -3783 -3538
rect -3786 -3544 -3783 -3541
rect -3786 -3547 -3765 -3544
rect -3756 -3560 -3753 -3550
rect -3819 -3563 -3753 -3560
rect -3819 -3581 -3816 -3563
rect -5979 -3604 -5708 -3599
rect -5703 -3604 -4923 -3599
rect -6097 -3655 -6094 -3649
rect -6097 -3658 -6060 -3655
rect -6063 -3661 -6060 -3658
rect -6063 -3664 -6042 -3661
rect -4652 -3666 -4293 -3661
rect -4279 -3665 -3829 -3660
rect -3816 -3666 -3813 -3660
rect -6033 -3677 -6030 -3667
rect -3816 -3669 -3779 -3666
rect -3782 -3672 -3779 -3669
rect -6096 -3680 -6030 -3677
rect -6096 -3698 -6093 -3680
rect -3782 -3675 -3761 -3672
rect -3752 -3688 -3749 -3678
rect -7704 -3704 -6430 -3699
rect -6425 -3704 -6185 -3699
rect -3815 -3691 -3749 -3688
rect -3815 -3709 -3812 -3691
rect -5877 -3783 -5087 -3778
rect -6094 -3799 -6091 -3793
rect -6094 -3802 -6057 -3799
rect -6060 -3805 -6057 -3802
rect -6060 -3808 -6039 -3805
rect -4535 -3809 -4294 -3804
rect -4280 -3808 -3828 -3803
rect -3815 -3809 -3812 -3803
rect -6030 -3821 -6027 -3811
rect -3815 -3812 -3778 -3809
rect -3781 -3815 -3778 -3812
rect -6093 -3824 -6027 -3821
rect -6093 -3842 -6090 -3824
rect -3781 -3818 -3760 -3815
rect -3751 -3831 -3748 -3821
rect -5976 -3838 -5616 -3833
rect -5611 -3838 -4749 -3833
rect -3814 -3834 -3748 -3831
rect -7838 -3848 -6485 -3843
rect -6480 -3848 -6183 -3843
rect -3814 -3852 -3811 -3834
rect -5980 -3869 -5487 -3864
rect -5482 -3869 -4625 -3864
rect -6098 -3947 -6095 -3941
rect -6098 -3950 -6061 -3947
rect -6064 -3953 -6061 -3950
rect -6064 -3956 -6043 -3953
rect -6034 -3969 -6031 -3959
rect -4393 -3961 -4294 -3956
rect -4280 -3960 -3610 -3955
rect -6097 -3972 -6031 -3969
rect -6097 -3990 -6094 -3972
rect -7980 -3996 -6546 -3991
rect -6541 -3996 -6179 -3991
rect -5955 -4032 -5327 -4027
rect -5322 -4032 -4485 -4027
rect -6073 -4163 -6070 -4157
rect -6073 -4166 -6036 -4163
rect -6039 -4169 -6036 -4166
rect -6039 -4172 -6018 -4169
rect -6009 -4185 -6006 -4175
rect -6072 -4188 -6006 -4185
rect -6072 -4206 -6069 -4188
rect -8122 -4212 -6597 -4207
rect -6592 -4212 -6154 -4207
rect -5984 -4407 -4914 -4402
rect -6368 -4413 -6213 -4409
rect -6383 -4418 -6221 -4417
rect -6383 -4422 -6219 -4418
rect -6219 -4425 -6213 -4423
rect -5991 -4440 -4740 -4435
rect -5972 -4511 -4616 -4506
rect -6146 -4522 -6121 -4518
rect -6412 -4523 -6121 -4522
rect -6412 -4526 -6140 -4523
rect -6425 -4534 -6121 -4530
rect -6425 -4535 -6114 -4534
rect -5951 -4610 -4477 -4605
rect -6158 -4647 -6136 -4646
rect -6465 -4651 -6136 -4647
rect -6480 -4660 -6134 -4655
rect -6128 -4660 -6127 -4655
rect -5932 -4669 -4398 -4664
rect -6156 -4769 -6128 -4765
rect -6524 -4771 -6128 -4769
rect -6122 -4771 -6121 -4767
rect -6524 -4772 -6121 -4771
rect -6524 -4773 -6154 -4772
rect -6541 -4781 -6128 -4777
rect -6122 -4781 -6121 -4777
rect -6541 -4782 -6121 -4781
rect -6154 -4910 -6126 -4906
rect -6580 -4912 -6126 -4910
rect -6120 -4912 -6119 -4908
rect -6580 -4913 -6119 -4912
rect -6580 -4914 -6152 -4913
rect -6592 -4922 -6126 -4918
rect -6120 -4922 -6119 -4918
rect -6592 -4923 -6119 -4922
rect -5241 -4927 -5231 -4922
rect -5081 -4927 -5078 -4922
<< m3contact >>
rect -6373 -3477 -6368 -3472
rect -6388 -3532 -6383 -3527
rect -6417 -3650 -6412 -3645
rect -6430 -3704 -6425 -3699
rect -6470 -3794 -6465 -3789
rect -6485 -3848 -6480 -3843
rect -6529 -3942 -6524 -3937
rect -6546 -3996 -6541 -3991
rect -6585 -4158 -6580 -4153
rect -6597 -4212 -6592 -4207
rect -6470 -4651 -6465 -4646
rect -6485 -4660 -6480 -4655
rect -6529 -4773 -6524 -4768
rect -6546 -4782 -6541 -4777
rect -6585 -4914 -6580 -4909
rect -6597 -4923 -6592 -4918
<< m123contact >>
rect -3739 -3187 -3734 -3182
rect -3739 -3240 -3734 -3235
rect -3721 -3236 -3716 -3231
rect -3707 -3281 -3702 -3276
rect -3808 -3371 -3803 -3366
rect -3808 -3424 -3803 -3419
rect -3790 -3420 -3785 -3415
rect -6083 -3446 -6078 -3441
rect -3776 -3465 -3771 -3460
rect -6083 -3499 -6078 -3494
rect -6065 -3495 -6060 -3490
rect -3813 -3501 -3808 -3496
rect -6051 -3540 -6046 -3535
rect -3813 -3554 -3808 -3549
rect -3795 -3550 -3790 -3545
rect -3781 -3595 -3776 -3590
rect -6090 -3618 -6085 -3613
rect -3809 -3629 -3804 -3624
rect -6090 -3671 -6085 -3666
rect -6072 -3667 -6067 -3662
rect -3809 -3682 -3804 -3677
rect -3791 -3678 -3786 -3673
rect -6058 -3712 -6053 -3707
rect -3777 -3723 -3772 -3718
rect -6087 -3762 -6082 -3757
rect -3808 -3772 -3803 -3767
rect -6087 -3815 -6082 -3810
rect -6069 -3811 -6064 -3806
rect -3808 -3825 -3803 -3820
rect -3790 -3821 -3785 -3816
rect -6055 -3856 -6050 -3851
rect -3776 -3866 -3771 -3861
rect -6091 -3910 -6086 -3905
rect -6091 -3963 -6086 -3958
rect -6073 -3959 -6068 -3954
rect -6059 -4004 -6054 -3999
rect -6066 -4126 -6061 -4121
rect -6066 -4179 -6061 -4174
rect -6048 -4175 -6043 -4170
rect -6034 -4220 -6029 -4215
rect -6373 -4413 -6368 -4408
rect -6388 -4422 -6383 -4417
rect -6417 -4526 -6412 -4521
rect -6430 -4535 -6425 -4530
<< metal3 >>
rect -3739 -3235 -3736 -3187
rect -3716 -3236 -3704 -3233
rect -3707 -3276 -3704 -3236
rect -3808 -3419 -3805 -3371
rect -3785 -3420 -3773 -3417
rect -6470 -3789 -6465 -3788
rect -6529 -3937 -6524 -3936
rect -6597 -4918 -6592 -4212
rect -6585 -4909 -6580 -4158
rect -6546 -4777 -6541 -3996
rect -6529 -4768 -6524 -3942
rect -6485 -4655 -6480 -3848
rect -6470 -4646 -6465 -3794
rect -6430 -4530 -6425 -3704
rect -6417 -4521 -6412 -3650
rect -6388 -4417 -6383 -3532
rect -6373 -4408 -6368 -3477
rect -6083 -3494 -6080 -3446
rect -3776 -3460 -3773 -3420
rect -6060 -3495 -6048 -3492
rect -6051 -3535 -6048 -3495
rect -3813 -3549 -3810 -3501
rect -3790 -3550 -3778 -3547
rect -3781 -3590 -3778 -3550
rect -6090 -3666 -6087 -3618
rect -6067 -3667 -6055 -3664
rect -6058 -3707 -6055 -3667
rect -3809 -3677 -3806 -3629
rect -3786 -3678 -3774 -3675
rect -3777 -3718 -3774 -3678
rect -6087 -3810 -6084 -3762
rect -6064 -3811 -6052 -3808
rect -6055 -3851 -6052 -3811
rect -3808 -3820 -3805 -3772
rect -3785 -3821 -3773 -3818
rect -3776 -3861 -3773 -3821
rect -6091 -3958 -6088 -3910
rect -6068 -3959 -6056 -3956
rect -6059 -3999 -6056 -3959
rect -6066 -4174 -6063 -4126
rect -6043 -4175 -6031 -4172
rect -6034 -4215 -6031 -4175
rect -6470 -4652 -6465 -4651
<< labels >>
rlabel metal2 -3610 -3958 -3609 -3957 1 cout
rlabel metal1 -4294 -3994 -4290 -3990 1 gnd!
rlabel metal1 -4294 -3896 -4290 -3893 1 vdd!
rlabel metal1 -5958 -4033 -5958 -4031 1 prop_5
rlabel metal1 -3721 -3287 -3717 -3284 1 gnd
rlabel metal1 -3671 -3281 -3668 -3279 1 gnd
rlabel metal1 -3723 -3231 -3722 -3229 1 gnd
rlabel metal1 -3727 -3187 -3724 -3185 5 vdd
rlabel metal1 -3726 -3241 -3723 -3239 1 vdd
rlabel metal1 -3630 -3250 -3630 -3250 1 s1
rlabel m2contact -3788 -3269 -3788 -3269 1 prop_1
rlabel metal1 -3701 -3836 -3699 -3834 1 s5
rlabel metal1 -3817 -3854 -3815 -3854 1 prop_5
rlabel metal1 -3795 -3826 -3792 -3824 1 vdd
rlabel metal1 -3796 -3772 -3793 -3770 5 vdd
rlabel metal1 -3792 -3816 -3791 -3814 1 gnd
rlabel metal1 -3740 -3866 -3737 -3864 1 gnd
rlabel metal1 -3790 -3872 -3786 -3869 1 gnd
rlabel metal1 -4390 -4662 -4386 -4657 7 clock_car0
rlabel metal1 -6013 -4873 -6013 -4873 5 vdd
rlabel metal1 -6010 -4930 -6010 -4930 1 gnd
rlabel metal1 -6042 -4948 -6042 -4948 1 gnd
rlabel metal1 -6043 -4861 -6043 -4861 5 vdd
rlabel metal1 -4493 -3207 -4489 -3202 5 vdd!
rlabel metal2 -4504 -3295 -4499 -3289 1 clock_in
rlabel metal1 -4469 -4603 -4465 -4598 7 clock_car0
rlabel metal2 -4485 -4610 -4481 -4605 1 gen_4
rlabel metal1 -4477 -4491 -4473 -4486 1 pdr4
rlabel metal1 -4477 -4046 -4473 -4016 1 pdr4
rlabel metal2 -4500 -4032 -4485 -4027 1 prop_5
rlabel metal1 -4485 -3916 -4481 -3899 1 pdr5
rlabel metal1 -6053 -4180 -6050 -4178 1 vdd
rlabel metal1 -6054 -4126 -6051 -4124 5 vdd
rlabel metal1 -6050 -4170 -6049 -4168 1 gnd
rlabel metal1 -5998 -4220 -5995 -4218 1 gnd
rlabel metal1 -6048 -4226 -6044 -4223 1 gnd
rlabel metal1 -5997 -4768 -5997 -4768 1 gen_4
rlabel metal1 -6015 -4732 -6015 -4732 5 vdd
rlabel metal1 -6012 -4789 -6012 -4789 1 gnd
rlabel metal1 -6044 -4807 -6044 -4807 1 gnd
rlabel metal1 -6045 -4720 -6045 -4720 5 vdd
rlabel metal1 -5974 -4648 -5974 -4648 1 gen_3
rlabel metal1 -6017 -4612 -6017 -4612 5 vdd
rlabel metal1 -6014 -4669 -6014 -4669 1 gnd
rlabel metal1 -6046 -4687 -6046 -4687 1 gnd
rlabel metal1 -6047 -4600 -6047 -4600 5 vdd
rlabel metal1 -5992 -4520 -5992 -4520 1 gen_2
rlabel metal1 -6020 -4484 -6020 -4484 5 vdd
rlabel metal1 -6017 -4541 -6017 -4541 1 gnd
rlabel metal1 -6049 -4559 -6049 -4559 1 gnd
rlabel metal1 -6050 -4472 -6050 -4472 5 vdd
rlabel metal1 -5985 -4412 -5985 -4412 1 gen_1
rlabel metal1 -6021 -4375 -6021 -4375 5 vdd
rlabel metal1 -6018 -4432 -6018 -4432 1 gnd
rlabel metal1 -6050 -4450 -6050 -4450 1 gnd
rlabel metal1 -6051 -4363 -6051 -4363 5 vdd
rlabel metal1 -5070 -4920 -5066 -4916 1 gnd!
rlabel metal1 -5078 -4807 -5074 -4803 1 clock_car0
rlabel metal1 -4608 -4504 -4604 -4500 1 clock_car0
rlabel metal2 -4624 -4511 -4620 -4506 1 gen_3
rlabel metal1 -4616 -4392 -4612 -4387 1 pdr3
rlabel metal1 -4906 -4400 -4902 -4396 1 clock_car0
rlabel metal2 -4922 -4407 -4918 -4402 1 gen_1
rlabel metal1 -4914 -4288 -4910 -4283 1 pdr1
rlabel metal1 -4732 -4433 -4728 -4428 1 clock_car0
rlabel metal2 -4748 -4440 -4744 -4435 1 gen_2
rlabel metal1 -4740 -4321 -4736 -4316 1 pdr2
rlabel metal1 -5879 -3172 -5879 -3172 1 carry_0
rlabel metal1 -3943 -3454 -3943 -3454 1 prop_2
rlabel metal1 -3819 -3711 -3819 -3711 1 prop_4
rlabel metal1 -3701 -3692 -3701 -3692 1 s4
rlabel metal1 -3796 -3683 -3793 -3681 1 vdd
rlabel metal1 -3797 -3629 -3794 -3627 5 vdd
rlabel metal1 -3793 -3673 -3792 -3671 1 gnd
rlabel metal1 -3741 -3723 -3738 -3721 1 gnd
rlabel metal1 -3791 -3729 -3787 -3726 1 gnd
rlabel metal1 -3830 -3529 -3830 -3529 1 c2
rlabel metal1 -3795 -3601 -3791 -3598 1 gnd
rlabel metal1 -3745 -3595 -3742 -3593 1 gnd
rlabel metal1 -3797 -3545 -3796 -3543 1 gnd
rlabel metal1 -3801 -3501 -3798 -3499 5 vdd
rlabel metal1 -3800 -3555 -3797 -3553 1 vdd
rlabel metal1 -3823 -3584 -3823 -3584 1 prop_3
rlabel metal1 -3704 -3564 -3704 -3564 1 s3
rlabel metal1 -3699 -3435 -3699 -3435 7 s2
rlabel metal1 -3817 -3400 -3817 -3400 1 c1
rlabel metal1 -3795 -3425 -3792 -3423 1 vdd
rlabel metal1 -3796 -3371 -3793 -3369 5 vdd
rlabel metal1 -3792 -3415 -3791 -3413 1 gnd
rlabel metal1 -3740 -3465 -3737 -3463 1 gnd
rlabel metal1 -3790 -3471 -3786 -3468 1 gnd
rlabel metal1 -5982 -3878 -5982 -3878 1 prop_4
rlabel metal1 -6078 -3964 -6075 -3962 1 vdd
rlabel metal1 -6079 -3910 -6076 -3908 5 vdd
rlabel metal1 -6075 -3954 -6074 -3952 1 gnd
rlabel metal1 -6023 -4004 -6020 -4002 1 gnd
rlabel metal1 -6073 -4010 -6069 -4007 1 gnd
rlabel metal1 -5979 -3825 -5979 -3825 1 prop_3
rlabel metal1 -6074 -3816 -6071 -3814 1 vdd
rlabel metal1 -6075 -3762 -6072 -3760 5 vdd
rlabel metal1 -6071 -3806 -6070 -3804 1 gnd
rlabel metal1 -6019 -3856 -6016 -3854 1 gnd
rlabel metal1 -6069 -3862 -6065 -3859 1 gnd
rlabel metal1 -5982 -3680 -5982 -3680 1 prop_2
rlabel metal1 -6077 -3672 -6074 -3670 1 vdd
rlabel metal1 -6078 -3618 -6075 -3616 5 vdd
rlabel metal1 -6074 -3662 -6073 -3660 1 gnd
rlabel metal1 -6022 -3712 -6019 -3710 1 gnd
rlabel metal1 -6072 -3718 -6068 -3715 1 gnd
rlabel metal1 -5977 -3509 -5977 -3509 1 prop_1
rlabel metal1 -6070 -3500 -6067 -3498 1 vdd
rlabel metal1 -6071 -3446 -6068 -3444 5 vdd
rlabel metal1 -6067 -3490 -6066 -3488 1 gnd
rlabel metal1 -6015 -3540 -6012 -3538 1 gnd
rlabel metal1 -6065 -3546 -6061 -3543 1 gnd
rlabel metal1 -4285 -3809 -4282 -3804 1 c4
rlabel metal2 -4297 -3809 -4295 -3804 1 pdr4
rlabel metal1 -4294 -3842 -4290 -3838 1 gnd!
rlabel metal1 -4294 -3744 -4290 -3741 1 vdd!
rlabel metal2 -4657 -3666 -4655 -3661 1 pdr3
rlabel metal1 -4284 -3666 -4281 -3661 1 c3
rlabel metal1 -4293 -3699 -4289 -3695 1 gnd!
rlabel metal1 -4293 -3601 -4289 -3598 1 vdd!
rlabel metal1 -4293 -3471 -4289 -3467 1 vdd!
rlabel metal1 -4293 -3568 -4289 -3564 1 gnd!
rlabel metal2 -4296 -3535 -4294 -3530 1 pdr2
rlabel m2contact -4284 -3535 -4281 -3530 1 c2
rlabel metal2 -4997 -3404 -4995 -3399 1 pdr1
rlabel metal1 -4285 -3404 -4282 -3400 1 c1
rlabel metal1 -4294 -3437 -4290 -3433 1 gnd!
rlabel metal1 -4294 -3340 -4290 -3336 1 vdd!
rlabel metal1 -4617 -3862 -4613 -3858 1 pdr3
rlabel metal2 -4633 -3869 -4629 -3864 1 prop_4
rlabel metal1 -4625 -3749 -4621 -3745 1 pdr4
rlabel metal1 -4741 -3831 -4737 -3827 1 pdr2
rlabel metal2 -4757 -3838 -4753 -3833 1 prop_3
rlabel metal1 -4749 -3719 -4745 -3714 1 pdr3
rlabel metal1 -5087 -3664 -5083 -3659 1 prop1_car0
rlabel metal2 -5095 -3783 -5091 -3778 1 carry_0
rlabel metal1 -5079 -3776 -5075 -3771 1 clock_car0
rlabel metal1 -5087 -3508 -5083 -3503 1 prop1_car0
rlabel metal2 -5103 -3515 -5098 -3510 2 prop_1
rlabel metal1 -5095 -3396 -5091 -3391 1 pdr1
rlabel metal1 -4915 -3597 -4911 -3592 1 pdr1
rlabel metal2 -4931 -3604 -4926 -3599 1 prop_2
rlabel metal1 -4923 -3485 -4919 -3480 1 pdr2
rlabel metal1 -4633 -3204 -4629 -3199 5 vdd!
rlabel metal2 -4644 -3292 -4639 -3286 1 clock_in
rlabel metal1 -4625 -3283 -4621 -3279 1 pdr4
rlabel metal1 -4749 -3282 -4745 -3278 1 pdr3
rlabel metal2 -4768 -3291 -4762 -3285 1 clock_in
rlabel metal1 -4757 -3203 -4753 -3198 5 vdd!
rlabel metal1 -4931 -3203 -4927 -3198 5 vdd!
rlabel metal2 -4942 -3291 -4936 -3285 1 clock_in
rlabel metal1 -4923 -3282 -4919 -3278 1 pdr2
rlabel metal1 -5095 -3281 -5091 -3276 1 pdr1
rlabel metal2 -5114 -3290 -5108 -3284 2 clock_in
rlabel metal1 -5103 -3202 -5099 -3197 5 vdd!
rlabel metal1 -5228 -3045 -5225 -3041 1 clock_in
rlabel metal2 -5240 -3045 -5237 -3040 1 clk_org
rlabel metal1 -5237 -3078 -5233 -3074 1 gnd!
rlabel metal1 -5237 -2981 -5233 -2977 1 vdd!
rlabel metal1 -5996 -4910 -5994 -4908 1 gen_5
rlabel metal2 -4406 -4669 -4402 -4664 1 gen_5
rlabel metal2 -4297 -3961 -4295 -3956 1 pdr5
rlabel metal1 -4398 -4550 -4394 -4545 1 pdr5
rlabel metal1 -4485 -3286 -4481 -3282 1 pdr5
rlabel metal2 -5086 -4927 -5081 -4922 1 clock_in
rlabel metal1 -5222 -4927 -5219 -4923 1 clock_in
rlabel metal2 -5234 -4927 -5231 -4922 1 clk_org
rlabel metal1 -5231 -4960 -5227 -4956 1 gnd!
rlabel metal1 -5231 -4863 -5227 -4859 1 vdd!
rlabel metal1 -3372 -3225 -3371 -3223 1 vdd!
rlabel metal1 -3372 -3271 -3371 -3269 1 gnd!
rlabel metal1 -3564 -3229 -3539 -3225 1 vdd!
rlabel metal1 -3564 -3267 -3539 -3264 1 gnd!
rlabel metal1 -3464 -3266 -3463 -3265 1 gnd!
rlabel metal1 -3469 -3227 -3468 -3226 1 vdd!
rlabel metal1 -3156 -3225 -3155 -3223 1 vdd!
rlabel metal1 -3156 -3271 -3155 -3269 1 gnd!
rlabel metal1 -3348 -3229 -3323 -3225 1 vdd!
rlabel metal1 -3348 -3267 -3323 -3264 1 gnd!
rlabel metal1 -3248 -3266 -3247 -3265 1 gnd!
rlabel metal1 -3253 -3227 -3252 -3226 1 vdd!
rlabel metal1 -3310 -3218 -3307 -3214 5 clock_org
rlabel metal1 -3312 -3275 -3309 -3271 1 clock_in
rlabel metal1 -3526 -3218 -3523 -3214 5 clock_org
rlabel metal1 -3528 -3275 -3524 -3271 1 clock_in
rlabel metal1 -3155 -3252 -3148 -3249 7 s1_final
rlabel metal1 -3377 -3409 -3376 -3407 1 vdd!
rlabel metal1 -3377 -3455 -3376 -3453 1 gnd!
rlabel metal1 -3569 -3413 -3544 -3409 1 vdd!
rlabel metal1 -3569 -3451 -3544 -3448 1 gnd!
rlabel metal1 -3469 -3450 -3468 -3449 1 gnd!
rlabel metal1 -3474 -3411 -3473 -3410 1 vdd!
rlabel metal1 -3161 -3409 -3160 -3407 1 vdd!
rlabel metal1 -3161 -3455 -3160 -3453 1 gnd!
rlabel metal1 -3353 -3413 -3328 -3409 1 vdd!
rlabel metal1 -3353 -3451 -3328 -3448 1 gnd!
rlabel metal1 -3253 -3450 -3252 -3449 1 gnd!
rlabel metal1 -3258 -3411 -3257 -3410 1 vdd!
rlabel metal1 -3315 -3402 -3312 -3398 5 clock_org
rlabel metal1 -3317 -3459 -3314 -3455 1 clock_in
rlabel metal1 -3531 -3402 -3528 -3398 5 clock_org
rlabel metal1 -3533 -3459 -3529 -3455 1 clock_in
rlabel metal1 -3160 -3436 -3153 -3433 1 s2_final
rlabel metal1 -3404 -3463 -3403 -3459 1 clock_org
rlabel metal1 -3405 -3398 -3404 -3396 1 clock_in
rlabel metal1 -3189 -3398 -3188 -3396 1 clock_org
rlabel metal1 -3188 -3463 -3187 -3459 1 clock_in
rlabel metal1 -3183 -3279 -3182 -3275 1 clock_in
rlabel metal1 -3184 -3214 -3183 -3212 1 clock_org
rlabel metal1 -3399 -3279 -3398 -3275 1 clock_org
rlabel metal1 -3400 -3214 -3399 -3212 1 clock_in
rlabel metal1 -3357 -3252 -3355 -3250 1 X1
rlabel metal1 -3363 -3436 -3360 -3434 1 X2
rlabel metal1 -3380 -3540 -3379 -3538 1 vdd!
rlabel metal1 -3380 -3586 -3379 -3584 1 gnd!
rlabel metal1 -3572 -3544 -3547 -3540 1 vdd!
rlabel metal1 -3572 -3582 -3547 -3579 1 gnd!
rlabel metal1 -3472 -3581 -3471 -3580 1 gnd!
rlabel metal1 -3477 -3542 -3476 -3541 1 vdd!
rlabel metal1 -3164 -3540 -3163 -3538 1 vdd!
rlabel metal1 -3164 -3586 -3163 -3584 1 gnd!
rlabel metal1 -3356 -3544 -3331 -3540 1 vdd!
rlabel metal1 -3356 -3582 -3331 -3579 1 gnd!
rlabel metal1 -3256 -3581 -3255 -3580 1 gnd!
rlabel metal1 -3261 -3542 -3260 -3541 1 vdd!
rlabel metal1 -3318 -3533 -3315 -3529 5 clock_org
rlabel metal1 -3320 -3590 -3317 -3586 1 clock_in
rlabel metal1 -3534 -3533 -3531 -3529 5 clock_org
rlabel metal1 -3536 -3590 -3532 -3586 1 clock_in
rlabel metal1 -3407 -3594 -3406 -3590 1 clock_org
rlabel metal1 -3408 -3529 -3407 -3527 1 clock_in
rlabel metal1 -3192 -3529 -3191 -3527 1 clock_org
rlabel metal1 -3191 -3594 -3190 -3590 1 clock_in
rlabel metal1 -3366 -3568 -3363 -3565 1 X3
rlabel metal1 -3163 -3567 -3156 -3564 1 s3_final
rlabel metal1 -3393 -3670 -3392 -3668 1 vdd!
rlabel metal1 -3393 -3716 -3392 -3714 1 gnd!
rlabel metal1 -3585 -3674 -3560 -3670 1 vdd!
rlabel metal1 -3585 -3712 -3560 -3709 1 gnd!
rlabel metal1 -3485 -3711 -3484 -3710 1 gnd!
rlabel metal1 -3490 -3672 -3489 -3671 1 vdd!
rlabel metal1 -3177 -3670 -3176 -3668 1 vdd!
rlabel metal1 -3177 -3716 -3176 -3714 1 gnd!
rlabel metal1 -3369 -3674 -3344 -3670 1 vdd!
rlabel metal1 -3369 -3712 -3344 -3709 1 gnd!
rlabel metal1 -3269 -3711 -3268 -3710 1 gnd!
rlabel metal1 -3274 -3672 -3273 -3671 1 vdd!
rlabel metal1 -3331 -3663 -3328 -3659 5 clock_org
rlabel metal1 -3333 -3720 -3330 -3716 1 clock_in
rlabel metal1 -3547 -3663 -3544 -3659 5 clock_org
rlabel metal1 -3549 -3720 -3545 -3716 1 clock_in
rlabel metal1 -3420 -3724 -3419 -3720 1 clock_org
rlabel metal1 -3421 -3659 -3420 -3657 1 clock_in
rlabel metal1 -3205 -3659 -3204 -3657 1 clock_org
rlabel metal1 -3204 -3724 -3203 -3720 1 clock_in
rlabel metal1 -3392 -3813 -3391 -3811 1 vdd!
rlabel metal1 -3392 -3859 -3391 -3857 1 gnd!
rlabel metal1 -3584 -3817 -3559 -3813 1 vdd!
rlabel metal1 -3584 -3855 -3559 -3852 1 gnd!
rlabel metal1 -3484 -3854 -3483 -3853 1 gnd!
rlabel metal1 -3489 -3815 -3488 -3814 1 vdd!
rlabel metal1 -3176 -3813 -3175 -3811 1 vdd!
rlabel metal1 -3176 -3859 -3175 -3857 1 gnd!
rlabel metal1 -3368 -3817 -3343 -3813 1 vdd!
rlabel metal1 -3368 -3855 -3343 -3852 1 gnd!
rlabel metal1 -3268 -3854 -3267 -3853 1 gnd!
rlabel metal1 -3273 -3815 -3272 -3814 1 vdd!
rlabel metal1 -3330 -3806 -3327 -3802 5 clock_org
rlabel metal1 -3332 -3863 -3329 -3859 1 clock_in
rlabel metal1 -3546 -3806 -3543 -3802 5 clock_org
rlabel metal1 -3548 -3863 -3544 -3859 1 clock_in
rlabel metal1 -3419 -3867 -3418 -3863 1 clock_org
rlabel metal1 -3420 -3802 -3419 -3800 1 clock_in
rlabel metal1 -3204 -3802 -3203 -3800 1 clock_org
rlabel metal1 -3203 -3867 -3202 -3863 1 clock_in
rlabel metal1 -3407 -3931 -3406 -3929 1 vdd!
rlabel metal1 -3407 -3977 -3406 -3975 1 gnd!
rlabel metal1 -3599 -3935 -3574 -3931 1 vdd!
rlabel metal1 -3599 -3973 -3574 -3970 1 gnd!
rlabel metal1 -3499 -3972 -3498 -3971 1 gnd!
rlabel metal1 -3504 -3933 -3503 -3932 1 vdd!
rlabel metal1 -3191 -3931 -3190 -3929 1 vdd!
rlabel metal1 -3191 -3977 -3190 -3975 1 gnd!
rlabel metal1 -3383 -3935 -3358 -3931 1 vdd!
rlabel metal1 -3383 -3973 -3358 -3970 1 gnd!
rlabel metal1 -3283 -3972 -3282 -3971 1 gnd!
rlabel metal1 -3288 -3933 -3287 -3932 1 vdd!
rlabel metal1 -3345 -3924 -3342 -3920 5 clock_org
rlabel metal1 -3347 -3981 -3344 -3977 1 clock_in
rlabel metal1 -3561 -3924 -3558 -3920 5 clock_org
rlabel metal1 -3563 -3981 -3559 -3977 1 clock_in
rlabel metal1 -3434 -3985 -3433 -3981 1 clock_org
rlabel metal1 -3435 -3920 -3434 -3918 1 clock_in
rlabel metal1 -3219 -3920 -3218 -3918 1 clock_org
rlabel metal1 -3218 -3985 -3217 -3981 1 clock_in
rlabel metal1 -3176 -3697 -3169 -3694 1 s4_final
rlabel metal1 -3175 -3840 -3168 -3837 1 s5_final
rlabel metal1 -3190 -3958 -3183 -3955 1 cout_final
rlabel metal1 -3393 -3959 -3390 -3956 1 Xc
rlabel metal1 -3378 -3841 -3375 -3838 1 X5
rlabel metal1 -3379 -3698 -3376 -3695 1 X4
rlabel metal1 -7810 -3033 -7808 -3032 3 vdd!
rlabel metal1 -7856 -3033 -7854 -3032 3 gnd!
rlabel metal1 -7799 -3005 -7797 -3004 3 clock_org
rlabel metal1 -7864 -3006 -7860 -3005 3 clock_in
rlabel metal1 -7814 -2649 -7810 -2624 3 vdd!
rlabel metal1 -7852 -2649 -7849 -2624 3 gnd!
rlabel metal1 -7864 -2790 -7860 -2789 3 clock_org
rlabel metal1 -7860 -2879 -7856 -2876 3 clock_in
rlabel metal1 -7860 -2664 -7856 -2660 3 clock_in
rlabel metal1 -7799 -2789 -7797 -2788 3 clock_in
rlabel metal1 -7803 -2665 -7799 -2662 7 clock_org
rlabel metal1 -7803 -2881 -7799 -2878 7 clock_org
rlabel metal1 -7812 -2936 -7811 -2935 3 vdd!
rlabel metal1 -7851 -2941 -7850 -2940 3 gnd!
rlabel metal1 -7852 -2865 -7849 -2840 3 gnd!
rlabel metal1 -7814 -2865 -7810 -2840 3 vdd!
rlabel metal1 -7812 -2720 -7811 -2719 3 vdd!
rlabel metal1 -7851 -2725 -7850 -2724 3 gnd!
rlabel metal1 -7856 -2817 -7854 -2816 3 gnd!
rlabel metal1 -7810 -2817 -7808 -2816 3 vdd!
rlabel metal1 -7676 -3026 -7674 -3025 3 vdd!
rlabel metal1 -7722 -3026 -7720 -3025 3 gnd!
rlabel metal1 -7665 -2998 -7663 -2997 3 clock_org
rlabel metal1 -7730 -2999 -7726 -2998 3 clock_in
rlabel metal1 -7680 -2642 -7676 -2617 3 vdd!
rlabel metal1 -7718 -2642 -7715 -2617 3 gnd!
rlabel metal1 -7730 -2783 -7726 -2782 3 clock_org
rlabel metal1 -7726 -2872 -7722 -2869 3 clock_in
rlabel metal1 -7726 -2657 -7722 -2653 3 clock_in
rlabel metal1 -7665 -2782 -7663 -2781 3 clock_in
rlabel metal1 -7669 -2658 -7665 -2655 7 clock_org
rlabel metal1 -7669 -2874 -7665 -2871 7 clock_org
rlabel metal1 -7678 -2929 -7677 -2928 3 vdd!
rlabel metal1 -7717 -2934 -7716 -2933 3 gnd!
rlabel metal1 -7718 -2858 -7715 -2833 3 gnd!
rlabel metal1 -7680 -2858 -7676 -2833 3 vdd!
rlabel metal1 -7678 -2713 -7677 -2712 3 vdd!
rlabel metal1 -7717 -2718 -7716 -2717 3 gnd!
rlabel metal1 -7722 -2810 -7720 -2809 3 gnd!
rlabel metal1 -7676 -2810 -7674 -2809 3 vdd!
rlabel metal1 -7541 -3032 -7539 -3031 3 vdd!
rlabel metal1 -7587 -3032 -7585 -3031 3 gnd!
rlabel metal1 -7530 -3004 -7528 -3003 3 clock_org
rlabel metal1 -7595 -3005 -7591 -3004 3 clock_in
rlabel metal1 -7545 -2648 -7541 -2623 3 vdd!
rlabel metal1 -7583 -2648 -7580 -2623 3 gnd!
rlabel metal1 -7595 -2789 -7591 -2788 3 clock_org
rlabel metal1 -7591 -2878 -7587 -2875 3 clock_in
rlabel metal1 -7591 -2663 -7587 -2659 3 clock_in
rlabel metal1 -7530 -2788 -7528 -2787 3 clock_in
rlabel metal1 -7534 -2664 -7530 -2661 7 clock_org
rlabel metal1 -7534 -2880 -7530 -2877 7 clock_org
rlabel metal1 -7543 -2935 -7542 -2934 3 vdd!
rlabel metal1 -7582 -2940 -7581 -2939 3 gnd!
rlabel metal1 -7583 -2864 -7580 -2839 3 gnd!
rlabel metal1 -7545 -2864 -7541 -2839 3 vdd!
rlabel metal1 -7543 -2719 -7542 -2718 3 vdd!
rlabel metal1 -7582 -2724 -7581 -2723 3 gnd!
rlabel metal1 -7587 -2816 -7585 -2815 3 gnd!
rlabel metal1 -7541 -2816 -7539 -2815 3 vdd!
rlabel metal1 -7421 -3031 -7419 -3030 3 vdd!
rlabel metal1 -7467 -3031 -7465 -3030 3 gnd!
rlabel metal1 -7410 -3003 -7408 -3002 3 clock_org
rlabel metal1 -7475 -3004 -7471 -3003 3 clock_in
rlabel metal1 -7425 -2647 -7421 -2622 3 vdd!
rlabel metal1 -7463 -2647 -7460 -2622 3 gnd!
rlabel metal1 -7475 -2788 -7471 -2787 3 clock_org
rlabel metal1 -7471 -2877 -7467 -2874 3 clock_in
rlabel metal1 -7471 -2662 -7467 -2658 3 clock_in
rlabel metal1 -7410 -2787 -7408 -2786 3 clock_in
rlabel metal1 -7414 -2663 -7410 -2660 7 clock_org
rlabel metal1 -7414 -2879 -7410 -2876 7 clock_org
rlabel metal1 -7423 -2934 -7422 -2933 3 vdd!
rlabel metal1 -7462 -2939 -7461 -2938 3 gnd!
rlabel metal1 -7463 -2863 -7460 -2838 3 gnd!
rlabel metal1 -7425 -2863 -7421 -2838 3 vdd!
rlabel metal1 -7423 -2718 -7422 -2717 3 vdd!
rlabel metal1 -7462 -2723 -7461 -2722 3 gnd!
rlabel metal1 -7467 -2815 -7465 -2814 3 gnd!
rlabel metal1 -7421 -2815 -7419 -2814 3 vdd!
rlabel metal1 -7301 -3031 -7299 -3030 3 vdd!
rlabel metal1 -7347 -3031 -7345 -3030 3 gnd!
rlabel metal1 -7290 -3003 -7288 -3002 3 clock_org
rlabel metal1 -7355 -3004 -7351 -3003 3 clock_in
rlabel metal1 -7305 -2647 -7301 -2622 3 vdd!
rlabel metal1 -7343 -2647 -7340 -2622 3 gnd!
rlabel metal1 -7355 -2788 -7351 -2787 3 clock_org
rlabel metal1 -7351 -2877 -7347 -2874 3 clock_in
rlabel metal1 -7351 -2662 -7347 -2658 3 clock_in
rlabel metal1 -7290 -2787 -7288 -2786 3 clock_in
rlabel metal1 -7294 -2663 -7290 -2660 7 clock_org
rlabel metal1 -7294 -2879 -7290 -2876 7 clock_org
rlabel metal1 -7303 -2934 -7302 -2933 3 vdd!
rlabel metal1 -7342 -2939 -7341 -2938 3 gnd!
rlabel metal1 -7343 -2863 -7340 -2838 3 gnd!
rlabel metal1 -7305 -2863 -7301 -2838 3 vdd!
rlabel metal1 -7303 -2718 -7302 -2717 3 vdd!
rlabel metal1 -7342 -2723 -7341 -2722 3 gnd!
rlabel metal1 -7347 -2815 -7345 -2814 3 gnd!
rlabel metal1 -7301 -2815 -7299 -2814 3 vdd!
rlabel metal1 -7176 -3030 -7174 -3029 3 vdd!
rlabel metal1 -7222 -3030 -7220 -3029 3 gnd!
rlabel metal1 -7165 -3002 -7163 -3001 3 clock_org
rlabel metal1 -7230 -3003 -7226 -3002 3 clock_in
rlabel metal1 -7180 -2646 -7176 -2621 3 vdd!
rlabel metal1 -7218 -2646 -7215 -2621 3 gnd!
rlabel metal1 -7230 -2787 -7226 -2786 3 clock_org
rlabel metal1 -7226 -2876 -7222 -2873 3 clock_in
rlabel metal1 -7226 -2661 -7222 -2657 3 clock_in
rlabel metal1 -7165 -2786 -7163 -2785 3 clock_in
rlabel metal1 -7169 -2662 -7165 -2659 7 clock_org
rlabel metal1 -7169 -2878 -7165 -2875 7 clock_org
rlabel metal1 -7178 -2933 -7177 -2932 3 vdd!
rlabel metal1 -7217 -2938 -7216 -2937 3 gnd!
rlabel metal1 -7218 -2862 -7215 -2837 3 gnd!
rlabel metal1 -7180 -2862 -7176 -2837 3 vdd!
rlabel metal1 -7178 -2717 -7177 -2716 3 vdd!
rlabel metal1 -7217 -2722 -7216 -2721 3 gnd!
rlabel metal1 -7222 -2814 -7220 -2813 3 gnd!
rlabel metal1 -7176 -2814 -7174 -2813 3 vdd!
rlabel metal1 -7058 -3030 -7056 -3029 3 vdd!
rlabel metal1 -7104 -3030 -7102 -3029 3 gnd!
rlabel metal1 -7047 -3002 -7045 -3001 3 clock_org
rlabel metal1 -7112 -3003 -7108 -3002 3 clock_in
rlabel metal1 -7062 -2646 -7058 -2621 3 vdd!
rlabel metal1 -7100 -2646 -7097 -2621 3 gnd!
rlabel metal1 -7112 -2787 -7108 -2786 3 clock_org
rlabel metal1 -7108 -2876 -7104 -2873 3 clock_in
rlabel metal1 -7108 -2661 -7104 -2657 3 clock_in
rlabel metal1 -7047 -2786 -7045 -2785 3 clock_in
rlabel metal1 -7051 -2662 -7047 -2659 7 clock_org
rlabel metal1 -7051 -2878 -7047 -2875 7 clock_org
rlabel metal1 -7060 -2933 -7059 -2932 3 vdd!
rlabel metal1 -7099 -2938 -7098 -2937 3 gnd!
rlabel metal1 -7100 -2862 -7097 -2837 3 gnd!
rlabel metal1 -7062 -2862 -7058 -2837 3 vdd!
rlabel metal1 -7060 -2717 -7059 -2716 3 vdd!
rlabel metal1 -7099 -2722 -7098 -2721 3 gnd!
rlabel metal1 -7104 -2814 -7102 -2813 3 gnd!
rlabel metal1 -7058 -2814 -7056 -2813 3 vdd!
rlabel metal1 -6939 -3028 -6937 -3027 3 vdd!
rlabel metal1 -6985 -3028 -6983 -3027 3 gnd!
rlabel metal1 -6928 -3000 -6926 -2999 3 clock_org
rlabel metal1 -6993 -3001 -6989 -3000 3 clock_in
rlabel metal1 -6943 -2644 -6939 -2619 3 vdd!
rlabel metal1 -6981 -2644 -6978 -2619 3 gnd!
rlabel metal1 -6993 -2785 -6989 -2784 3 clock_org
rlabel metal1 -6989 -2874 -6985 -2871 3 clock_in
rlabel metal1 -6989 -2659 -6985 -2655 3 clock_in
rlabel metal1 -6967 -2613 -6963 -2608 5 q_a1
rlabel metal1 -6928 -2784 -6926 -2783 3 clock_in
rlabel metal1 -6932 -2660 -6928 -2657 7 clock_org
rlabel metal1 -6932 -2876 -6928 -2873 7 clock_org
rlabel metal1 -6941 -2931 -6940 -2930 3 vdd!
rlabel metal1 -6980 -2936 -6979 -2935 3 gnd!
rlabel metal1 -6981 -2860 -6978 -2835 3 gnd!
rlabel metal1 -6943 -2860 -6939 -2835 3 vdd!
rlabel metal1 -6941 -2715 -6940 -2714 3 vdd!
rlabel metal1 -6980 -2720 -6979 -2719 3 gnd!
rlabel metal1 -6985 -2812 -6983 -2811 3 gnd!
rlabel metal1 -6939 -2812 -6937 -2811 3 vdd!
rlabel metal1 -7086 -2615 -7082 -2610 1 q_a2
rlabel metal1 -7204 -2615 -7200 -2610 1 q_a3
rlabel metal1 -7329 -2616 -7325 -2611 1 q_a4
rlabel metal1 -7449 -2616 -7445 -2611 1 q_a5
rlabel metal1 -7569 -2617 -7565 -2612 1 q_b1
rlabel metal1 -7704 -2611 -7700 -2606 1 q_b2
rlabel metal1 -7838 -2618 -7834 -2613 1 q_b3
rlabel metal1 -8094 -3032 -8092 -3031 3 vdd!
rlabel metal1 -8140 -3032 -8138 -3031 3 gnd!
rlabel metal1 -8083 -3004 -8081 -3003 3 clock_org
rlabel metal1 -8148 -3005 -8144 -3004 3 clock_in
rlabel metal1 -8098 -2648 -8094 -2623 3 vdd!
rlabel metal1 -8136 -2648 -8133 -2623 3 gnd!
rlabel metal1 -8148 -2789 -8144 -2788 3 clock_org
rlabel metal1 -8144 -2878 -8140 -2875 3 clock_in
rlabel metal1 -8144 -2663 -8140 -2659 3 clock_in
rlabel metal1 -8083 -2788 -8081 -2787 3 clock_in
rlabel metal1 -8087 -2664 -8083 -2661 7 clock_org
rlabel metal1 -8087 -2880 -8083 -2877 7 clock_org
rlabel metal1 -8096 -2935 -8095 -2934 3 vdd!
rlabel metal1 -8135 -2940 -8134 -2939 3 gnd!
rlabel metal1 -8136 -2864 -8133 -2839 3 gnd!
rlabel metal1 -8098 -2864 -8094 -2839 3 vdd!
rlabel metal1 -8096 -2719 -8095 -2718 3 vdd!
rlabel metal1 -8135 -2724 -8134 -2723 3 gnd!
rlabel metal1 -8140 -2816 -8138 -2815 3 gnd!
rlabel metal1 -8094 -2816 -8092 -2815 3 vdd!
rlabel metal1 -7952 -3035 -7950 -3034 3 vdd!
rlabel metal1 -7998 -3035 -7996 -3034 3 gnd!
rlabel metal1 -7941 -3007 -7939 -3006 3 clock_org
rlabel metal1 -8006 -3008 -8002 -3007 3 clock_in
rlabel metal1 -7956 -2651 -7952 -2626 3 vdd!
rlabel metal1 -7994 -2651 -7991 -2626 3 gnd!
rlabel metal1 -8006 -2792 -8002 -2791 3 clock_org
rlabel metal1 -8002 -2881 -7998 -2878 3 clock_in
rlabel metal1 -8002 -2666 -7998 -2662 3 clock_in
rlabel metal1 -7941 -2791 -7939 -2790 3 clock_in
rlabel metal1 -7945 -2667 -7941 -2664 7 clock_org
rlabel metal1 -7945 -2883 -7941 -2880 7 clock_org
rlabel metal1 -7954 -2938 -7953 -2937 3 vdd!
rlabel metal1 -7993 -2943 -7992 -2942 3 gnd!
rlabel metal1 -7994 -2867 -7991 -2842 3 gnd!
rlabel metal1 -7956 -2867 -7952 -2842 3 vdd!
rlabel metal1 -7954 -2722 -7953 -2721 3 vdd!
rlabel metal1 -7993 -2727 -7992 -2726 3 gnd!
rlabel metal1 -7998 -2819 -7996 -2818 3 gnd!
rlabel metal1 -7952 -2819 -7950 -2818 3 vdd!
rlabel metal1 -7980 -2620 -7976 -2615 1 q_b4
rlabel metal1 -8122 -2617 -8118 -2612 1 q_b5
rlabel m2contact -6276 -3532 -6271 -3527 1 b1
rlabel metal1 -6270 -3476 -6268 -3473 1 a1
rlabel metal1 -6267 -3649 -6265 -3647 1 a2
rlabel m2contact -6184 -3702 -6182 -3700 1 b2
rlabel metal1 -6097 -3791 -6095 -3789 1 a3
rlabel metal1 -6097 -3845 -6095 -3843 1 b3
rlabel metal1 -6179 -3940 -6177 -3938 1 a4
rlabel m2contact -6179 -3993 -6177 -3991 1 b4
rlabel metal1 -6171 -4156 -6169 -4154 1 a5
rlabel m2contact -6154 -4212 -6149 -4207 1 b5
rlabel m2contact -6213 -4414 -6208 -4409 1 a1
rlabel m2contact -6120 -4523 -6117 -4520 1 a2
rlabel metal1 -6120 -4530 -6117 -4527 1 b2
rlabel m2contact -6215 -4420 -6214 -4419 1 b1
rlabel m2contact -6136 -4651 -6134 -4649 1 a3
rlabel m2contact -6132 -4657 -6130 -4655 1 b3
rlabel m2contact -6127 -4770 -6125 -4768 1 a4
rlabel metal1 -6127 -4776 -6125 -4774 1 b4
rlabel m2contact -6126 -4912 -6120 -4906 1 a5
rlabel metal1 -6126 -4922 -6120 -4916 1 b5
rlabel metal1 -6967 -2829 -6963 -2825 1 i1
rlabel metal1 -7086 -2831 -7082 -2827 1 i2
rlabel metal1 -7204 -2831 -7200 -2827 1 i3
rlabel metal1 -7329 -2832 -7325 -2828 1 i4
rlabel metal1 -7449 -2832 -7445 -2828 1 i5
rlabel metal1 -7569 -2833 -7565 -2829 1 i6
rlabel metal1 -7704 -2828 -7700 -2824 1 i7
rlabel metal1 -7838 -2834 -7834 -2830 1 i8
rlabel metal1 -7980 -2835 -7976 -2831 1 i9
rlabel metal1 -8122 -2833 -8118 -2829 1 i10
rlabel metal1 -6967 -3035 -6965 -3033 1 a1
rlabel metal1 -7085 -3037 -7083 -3035 1 a2
rlabel metal1 -7203 -3037 -7201 -3035 1 a3
rlabel metal1 -7329 -3037 -7327 -3035 1 a4
rlabel metal1 -7449 -3037 -7447 -3035 1 a5
rlabel metal1 -7568 -3036 -7566 -3034 1 b1
rlabel m2contact -7567 -3049 -7565 -3047 1 b1
rlabel m2contact -7703 -3039 -7701 -3037 1 b2
rlabel m2contact -7837 -3050 -7835 -3048 1 b3
rlabel m2contact -7978 -3052 -7976 -3050 1 b4
rlabel m2contact -8121 -3047 -8119 -3045 1 b5
<< end >>
