magic
tech scmos
timestamp 1763583544
<< nwell >>
rect -5243 -3036 -5219 -2984
rect -3739 -3211 -3715 -3187
rect -3700 -3197 -3666 -3191
rect -5109 -3273 -5085 -3211
rect -4937 -3274 -4913 -3212
rect -4763 -3274 -4739 -3212
rect -4639 -3275 -4615 -3213
rect -4499 -3278 -4475 -3216
rect -3700 -3227 -3638 -3197
rect -3672 -3233 -3638 -3227
rect -3739 -3266 -3715 -3242
rect -4300 -3395 -4276 -3343
rect -3808 -3395 -3784 -3371
rect -3769 -3381 -3735 -3375
rect -3769 -3411 -3707 -3381
rect -3741 -3417 -3707 -3411
rect -6083 -3470 -6059 -3446
rect -3808 -3450 -3784 -3426
rect -6044 -3456 -6010 -3450
rect -6044 -3486 -5982 -3456
rect -6016 -3492 -5982 -3486
rect -6083 -3525 -6059 -3501
rect -4299 -3526 -4275 -3474
rect -3813 -3525 -3789 -3501
rect -3774 -3511 -3740 -3505
rect -3774 -3541 -3712 -3511
rect -3746 -3547 -3712 -3541
rect -3813 -3580 -3789 -3556
rect -6090 -3642 -6066 -3618
rect -6051 -3628 -6017 -3622
rect -6051 -3658 -5989 -3628
rect -4299 -3657 -4275 -3605
rect -3809 -3653 -3785 -3629
rect -3770 -3639 -3736 -3633
rect -6023 -3664 -5989 -3658
rect -3770 -3669 -3708 -3639
rect -6090 -3697 -6066 -3673
rect -3742 -3675 -3708 -3669
rect -3809 -3708 -3785 -3684
rect -6087 -3786 -6063 -3762
rect -6048 -3772 -6014 -3766
rect -6048 -3802 -5986 -3772
rect -4300 -3800 -4276 -3748
rect -3808 -3796 -3784 -3772
rect -3769 -3782 -3735 -3776
rect -6020 -3808 -5986 -3802
rect -3769 -3812 -3707 -3782
rect -6087 -3841 -6063 -3817
rect -3741 -3818 -3707 -3812
rect -3808 -3851 -3784 -3827
rect -6091 -3934 -6067 -3910
rect -6052 -3920 -6018 -3914
rect -6052 -3950 -5990 -3920
rect -6024 -3956 -5990 -3950
rect -4300 -3952 -4276 -3900
rect -6091 -3989 -6067 -3965
rect -6066 -4150 -6042 -4126
rect -6027 -4136 -5993 -4130
rect -6027 -4166 -5965 -4136
rect -5999 -4172 -5965 -4166
rect -6066 -4205 -6042 -4181
rect -6067 -4401 -6031 -4361
rect -6025 -4408 -6001 -4368
rect -6066 -4510 -6030 -4470
rect -6024 -4517 -6000 -4477
rect -6063 -4638 -6027 -4598
rect -6021 -4645 -5997 -4605
rect -6061 -4758 -6025 -4718
rect -6019 -4765 -5995 -4725
rect -6059 -4899 -6023 -4859
rect -6017 -4906 -5993 -4866
rect -5237 -4918 -5213 -4866
<< ntransistor >>
rect -5232 -3068 -5230 -3048
rect -3728 -3225 -3726 -3219
rect -3689 -3274 -3687 -3262
rect -3679 -3274 -3677 -3262
rect -3661 -3274 -3659 -3262
rect -3651 -3274 -3649 -3262
rect -3728 -3280 -3726 -3274
rect -6072 -3484 -6070 -3478
rect -5090 -3499 -5088 -3399
rect -4289 -3427 -4287 -3407
rect -3797 -3409 -3795 -3403
rect -3758 -3458 -3756 -3446
rect -3748 -3458 -3746 -3446
rect -3730 -3458 -3728 -3446
rect -3720 -3458 -3718 -3446
rect -3797 -3464 -3795 -3458
rect -6033 -3533 -6031 -3521
rect -6023 -3533 -6021 -3521
rect -6005 -3533 -6003 -3521
rect -5995 -3533 -5993 -3521
rect -6072 -3539 -6070 -3533
rect -4918 -3588 -4916 -3488
rect -4288 -3558 -4286 -3538
rect -3802 -3539 -3800 -3533
rect -3763 -3588 -3761 -3576
rect -3753 -3588 -3751 -3576
rect -3735 -3588 -3733 -3576
rect -3725 -3588 -3723 -3576
rect -3802 -3594 -3800 -3588
rect -6079 -3656 -6077 -3650
rect -6040 -3705 -6038 -3693
rect -6030 -3705 -6028 -3693
rect -6012 -3705 -6010 -3693
rect -6002 -3705 -6000 -3693
rect -6079 -3711 -6077 -3705
rect -5082 -3767 -5080 -3667
rect -3798 -3667 -3796 -3661
rect -4288 -3689 -4286 -3669
rect -3759 -3716 -3757 -3704
rect -3749 -3716 -3747 -3704
rect -3731 -3716 -3729 -3704
rect -3721 -3716 -3719 -3704
rect -3798 -3722 -3796 -3716
rect -6076 -3800 -6074 -3794
rect -4744 -3822 -4742 -3722
rect -6037 -3849 -6035 -3837
rect -6027 -3849 -6025 -3837
rect -6009 -3849 -6007 -3837
rect -5999 -3849 -5997 -3837
rect -6076 -3855 -6074 -3849
rect -4620 -3853 -4618 -3753
rect -3797 -3810 -3795 -3804
rect -4289 -3832 -4287 -3812
rect -3758 -3859 -3756 -3847
rect -3748 -3859 -3746 -3847
rect -3730 -3859 -3728 -3847
rect -3720 -3859 -3718 -3847
rect -3797 -3865 -3795 -3859
rect -6080 -3948 -6078 -3942
rect -6041 -3997 -6039 -3985
rect -6031 -3997 -6029 -3985
rect -6013 -3997 -6011 -3985
rect -6003 -3997 -6001 -3985
rect -6080 -4003 -6078 -3997
rect -4480 -4016 -4478 -3916
rect -4289 -3984 -4287 -3964
rect -6055 -4164 -6053 -4158
rect -6016 -4213 -6014 -4201
rect -6006 -4213 -6004 -4201
rect -5988 -4213 -5986 -4201
rect -5978 -4213 -5976 -4201
rect -6055 -4219 -6053 -4213
rect -4909 -4391 -4907 -4291
rect -6056 -4444 -6054 -4424
rect -6045 -4444 -6043 -4424
rect -6014 -4426 -6012 -4416
rect -4735 -4424 -4733 -4324
rect -4611 -4495 -4609 -4395
rect -6055 -4553 -6053 -4533
rect -6044 -4553 -6042 -4533
rect -6013 -4535 -6011 -4525
rect -4472 -4594 -4470 -4494
rect -4393 -4653 -4391 -4553
rect -6052 -4681 -6050 -4661
rect -6041 -4681 -6039 -4661
rect -6010 -4663 -6008 -4653
rect -6050 -4801 -6048 -4781
rect -6039 -4801 -6037 -4781
rect -6008 -4783 -6006 -4773
rect -5073 -4911 -5071 -4811
rect -6048 -4942 -6046 -4922
rect -6037 -4942 -6035 -4922
rect -6006 -4924 -6004 -4914
rect -5226 -4950 -5224 -4930
<< ptransistor >>
rect -5232 -3030 -5230 -2990
rect -3728 -3205 -3726 -3193
rect -5098 -3267 -5096 -3217
rect -4926 -3268 -4924 -3218
rect -4752 -3268 -4750 -3218
rect -4628 -3269 -4626 -3219
rect -4488 -3272 -4486 -3222
rect -3689 -3221 -3687 -3197
rect -3679 -3221 -3677 -3197
rect -3661 -3227 -3659 -3203
rect -3651 -3227 -3649 -3203
rect -3728 -3260 -3726 -3248
rect -4289 -3389 -4287 -3349
rect -3797 -3389 -3795 -3377
rect -6072 -3464 -6070 -3452
rect -6033 -3480 -6031 -3456
rect -6023 -3480 -6021 -3456
rect -6005 -3486 -6003 -3462
rect -5995 -3486 -5993 -3462
rect -6072 -3519 -6070 -3507
rect -3758 -3405 -3756 -3381
rect -3748 -3405 -3746 -3381
rect -3730 -3411 -3728 -3387
rect -3720 -3411 -3718 -3387
rect -3797 -3444 -3795 -3432
rect -4288 -3520 -4286 -3480
rect -3802 -3519 -3800 -3507
rect -3763 -3535 -3761 -3511
rect -3753 -3535 -3751 -3511
rect -3735 -3541 -3733 -3517
rect -3725 -3541 -3723 -3517
rect -3802 -3574 -3800 -3562
rect -6079 -3636 -6077 -3624
rect -6040 -3652 -6038 -3628
rect -6030 -3652 -6028 -3628
rect -6012 -3658 -6010 -3634
rect -6002 -3658 -6000 -3634
rect -4288 -3651 -4286 -3611
rect -3798 -3647 -3796 -3635
rect -6079 -3691 -6077 -3679
rect -3759 -3663 -3757 -3639
rect -3749 -3663 -3747 -3639
rect -3731 -3669 -3729 -3645
rect -3721 -3669 -3719 -3645
rect -3798 -3702 -3796 -3690
rect -6076 -3780 -6074 -3768
rect -6037 -3796 -6035 -3772
rect -6027 -3796 -6025 -3772
rect -6009 -3802 -6007 -3778
rect -5999 -3802 -5997 -3778
rect -6076 -3835 -6074 -3823
rect -4289 -3794 -4287 -3754
rect -3797 -3790 -3795 -3778
rect -3758 -3806 -3756 -3782
rect -3748 -3806 -3746 -3782
rect -3730 -3812 -3728 -3788
rect -3720 -3812 -3718 -3788
rect -3797 -3845 -3795 -3833
rect -6080 -3928 -6078 -3916
rect -6041 -3944 -6039 -3920
rect -6031 -3944 -6029 -3920
rect -6013 -3950 -6011 -3926
rect -6003 -3950 -6001 -3926
rect -6080 -3983 -6078 -3971
rect -4289 -3946 -4287 -3906
rect -6055 -4144 -6053 -4132
rect -6016 -4160 -6014 -4136
rect -6006 -4160 -6004 -4136
rect -5988 -4166 -5986 -4142
rect -5978 -4166 -5976 -4142
rect -6055 -4199 -6053 -4187
rect -6056 -4395 -6054 -4375
rect -6045 -4395 -6043 -4375
rect -6014 -4402 -6012 -4382
rect -6055 -4504 -6053 -4484
rect -6044 -4504 -6042 -4484
rect -6013 -4511 -6011 -4491
rect -6052 -4632 -6050 -4612
rect -6041 -4632 -6039 -4612
rect -6010 -4639 -6008 -4619
rect -6050 -4752 -6048 -4732
rect -6039 -4752 -6037 -4732
rect -6008 -4759 -6006 -4739
rect -6048 -4893 -6046 -4873
rect -6037 -4893 -6035 -4873
rect -6006 -4900 -6004 -4880
rect -5226 -4912 -5224 -4872
<< ndiffusion >>
rect -5233 -3068 -5232 -3048
rect -5230 -3068 -5229 -3048
rect -3729 -3225 -3728 -3219
rect -3726 -3225 -3725 -3219
rect -3690 -3274 -3689 -3262
rect -3687 -3274 -3679 -3262
rect -3677 -3274 -3676 -3262
rect -3662 -3274 -3661 -3262
rect -3659 -3274 -3651 -3262
rect -3649 -3274 -3648 -3262
rect -3729 -3280 -3728 -3274
rect -3726 -3280 -3725 -3274
rect -6073 -3484 -6072 -3478
rect -6070 -3484 -6069 -3478
rect -5091 -3499 -5090 -3399
rect -5088 -3499 -5087 -3399
rect -4290 -3427 -4289 -3407
rect -4287 -3427 -4286 -3407
rect -3798 -3409 -3797 -3403
rect -3795 -3409 -3794 -3403
rect -3759 -3458 -3758 -3446
rect -3756 -3458 -3748 -3446
rect -3746 -3458 -3745 -3446
rect -3731 -3458 -3730 -3446
rect -3728 -3458 -3720 -3446
rect -3718 -3458 -3717 -3446
rect -3798 -3464 -3797 -3458
rect -3795 -3464 -3794 -3458
rect -6034 -3533 -6033 -3521
rect -6031 -3533 -6023 -3521
rect -6021 -3533 -6020 -3521
rect -6006 -3533 -6005 -3521
rect -6003 -3533 -5995 -3521
rect -5993 -3533 -5992 -3521
rect -6073 -3539 -6072 -3533
rect -6070 -3539 -6069 -3533
rect -4919 -3588 -4918 -3488
rect -4916 -3588 -4915 -3488
rect -4289 -3558 -4288 -3538
rect -4286 -3558 -4285 -3538
rect -3803 -3539 -3802 -3533
rect -3800 -3539 -3799 -3533
rect -3764 -3588 -3763 -3576
rect -3761 -3588 -3753 -3576
rect -3751 -3588 -3750 -3576
rect -3736 -3588 -3735 -3576
rect -3733 -3588 -3725 -3576
rect -3723 -3588 -3722 -3576
rect -3803 -3594 -3802 -3588
rect -3800 -3594 -3799 -3588
rect -6080 -3656 -6079 -3650
rect -6077 -3656 -6076 -3650
rect -6041 -3705 -6040 -3693
rect -6038 -3705 -6030 -3693
rect -6028 -3705 -6027 -3693
rect -6013 -3705 -6012 -3693
rect -6010 -3705 -6002 -3693
rect -6000 -3705 -5999 -3693
rect -6080 -3711 -6079 -3705
rect -6077 -3711 -6076 -3705
rect -5083 -3767 -5082 -3667
rect -5080 -3767 -5079 -3667
rect -3799 -3667 -3798 -3661
rect -3796 -3667 -3795 -3661
rect -4289 -3689 -4288 -3669
rect -4286 -3689 -4285 -3669
rect -3760 -3716 -3759 -3704
rect -3757 -3716 -3749 -3704
rect -3747 -3716 -3746 -3704
rect -3732 -3716 -3731 -3704
rect -3729 -3716 -3721 -3704
rect -3719 -3716 -3718 -3704
rect -3799 -3722 -3798 -3716
rect -3796 -3722 -3795 -3716
rect -6077 -3800 -6076 -3794
rect -6074 -3800 -6073 -3794
rect -4745 -3822 -4744 -3722
rect -4742 -3822 -4741 -3722
rect -6038 -3849 -6037 -3837
rect -6035 -3849 -6027 -3837
rect -6025 -3849 -6024 -3837
rect -6010 -3849 -6009 -3837
rect -6007 -3849 -5999 -3837
rect -5997 -3849 -5996 -3837
rect -6077 -3855 -6076 -3849
rect -6074 -3855 -6073 -3849
rect -4621 -3853 -4620 -3753
rect -4618 -3853 -4617 -3753
rect -3798 -3810 -3797 -3804
rect -3795 -3810 -3794 -3804
rect -4290 -3832 -4289 -3812
rect -4287 -3832 -4286 -3812
rect -3759 -3859 -3758 -3847
rect -3756 -3859 -3748 -3847
rect -3746 -3859 -3745 -3847
rect -3731 -3859 -3730 -3847
rect -3728 -3859 -3720 -3847
rect -3718 -3859 -3717 -3847
rect -3798 -3865 -3797 -3859
rect -3795 -3865 -3794 -3859
rect -6081 -3948 -6080 -3942
rect -6078 -3948 -6077 -3942
rect -6042 -3997 -6041 -3985
rect -6039 -3997 -6031 -3985
rect -6029 -3997 -6028 -3985
rect -6014 -3997 -6013 -3985
rect -6011 -3997 -6003 -3985
rect -6001 -3997 -6000 -3985
rect -6081 -4003 -6080 -3997
rect -6078 -4003 -6077 -3997
rect -4481 -4016 -4480 -3916
rect -4478 -4016 -4477 -3916
rect -4290 -3984 -4289 -3964
rect -4287 -3984 -4286 -3964
rect -6056 -4164 -6055 -4158
rect -6053 -4164 -6052 -4158
rect -6017 -4213 -6016 -4201
rect -6014 -4213 -6006 -4201
rect -6004 -4213 -6003 -4201
rect -5989 -4213 -5988 -4201
rect -5986 -4213 -5978 -4201
rect -5976 -4213 -5975 -4201
rect -6056 -4219 -6055 -4213
rect -6053 -4219 -6052 -4213
rect -4910 -4391 -4909 -4291
rect -4907 -4391 -4906 -4291
rect -6057 -4444 -6056 -4424
rect -6054 -4444 -6045 -4424
rect -6043 -4444 -6042 -4424
rect -6015 -4426 -6014 -4416
rect -6012 -4426 -6011 -4416
rect -4736 -4424 -4735 -4324
rect -4733 -4424 -4732 -4324
rect -4612 -4495 -4611 -4395
rect -4609 -4495 -4608 -4395
rect -6056 -4553 -6055 -4533
rect -6053 -4553 -6044 -4533
rect -6042 -4553 -6041 -4533
rect -6014 -4535 -6013 -4525
rect -6011 -4535 -6010 -4525
rect -4473 -4594 -4472 -4494
rect -4470 -4594 -4469 -4494
rect -4394 -4653 -4393 -4553
rect -4391 -4653 -4390 -4553
rect -6053 -4681 -6052 -4661
rect -6050 -4681 -6041 -4661
rect -6039 -4681 -6038 -4661
rect -6011 -4663 -6010 -4653
rect -6008 -4663 -6007 -4653
rect -6051 -4801 -6050 -4781
rect -6048 -4801 -6039 -4781
rect -6037 -4801 -6036 -4781
rect -6009 -4783 -6008 -4773
rect -6006 -4783 -6005 -4773
rect -5074 -4911 -5073 -4811
rect -5071 -4911 -5070 -4811
rect -6049 -4942 -6048 -4922
rect -6046 -4942 -6037 -4922
rect -6035 -4942 -6034 -4922
rect -6007 -4924 -6006 -4914
rect -6004 -4924 -6003 -4914
rect -5227 -4950 -5226 -4930
rect -5224 -4950 -5223 -4930
<< pdiffusion >>
rect -5233 -3030 -5232 -2990
rect -5230 -3030 -5229 -2990
rect -3729 -3205 -3728 -3193
rect -3726 -3205 -3725 -3193
rect -5099 -3267 -5098 -3217
rect -5096 -3267 -5095 -3217
rect -4927 -3268 -4926 -3218
rect -4924 -3268 -4923 -3218
rect -4753 -3268 -4752 -3218
rect -4750 -3268 -4749 -3218
rect -4629 -3269 -4628 -3219
rect -4626 -3269 -4625 -3219
rect -4489 -3272 -4488 -3222
rect -4486 -3272 -4485 -3222
rect -3690 -3221 -3689 -3197
rect -3687 -3221 -3685 -3197
rect -3681 -3221 -3679 -3197
rect -3677 -3221 -3676 -3197
rect -3662 -3227 -3661 -3203
rect -3659 -3227 -3657 -3203
rect -3653 -3227 -3651 -3203
rect -3649 -3227 -3648 -3203
rect -3729 -3260 -3728 -3248
rect -3726 -3260 -3725 -3248
rect -4290 -3389 -4289 -3349
rect -4287 -3389 -4286 -3349
rect -3798 -3389 -3797 -3377
rect -3795 -3389 -3794 -3377
rect -6073 -3464 -6072 -3452
rect -6070 -3464 -6069 -3452
rect -6034 -3480 -6033 -3456
rect -6031 -3480 -6029 -3456
rect -6025 -3480 -6023 -3456
rect -6021 -3480 -6020 -3456
rect -6006 -3486 -6005 -3462
rect -6003 -3486 -6001 -3462
rect -5997 -3486 -5995 -3462
rect -5993 -3486 -5992 -3462
rect -6073 -3519 -6072 -3507
rect -6070 -3519 -6069 -3507
rect -3759 -3405 -3758 -3381
rect -3756 -3405 -3754 -3381
rect -3750 -3405 -3748 -3381
rect -3746 -3405 -3745 -3381
rect -3731 -3411 -3730 -3387
rect -3728 -3411 -3726 -3387
rect -3722 -3411 -3720 -3387
rect -3718 -3411 -3717 -3387
rect -3798 -3444 -3797 -3432
rect -3795 -3444 -3794 -3432
rect -4289 -3520 -4288 -3480
rect -4286 -3520 -4285 -3480
rect -3803 -3519 -3802 -3507
rect -3800 -3519 -3799 -3507
rect -3764 -3535 -3763 -3511
rect -3761 -3535 -3759 -3511
rect -3755 -3535 -3753 -3511
rect -3751 -3535 -3750 -3511
rect -3736 -3541 -3735 -3517
rect -3733 -3541 -3731 -3517
rect -3727 -3541 -3725 -3517
rect -3723 -3541 -3722 -3517
rect -3803 -3574 -3802 -3562
rect -3800 -3574 -3799 -3562
rect -6080 -3636 -6079 -3624
rect -6077 -3636 -6076 -3624
rect -6041 -3652 -6040 -3628
rect -6038 -3652 -6036 -3628
rect -6032 -3652 -6030 -3628
rect -6028 -3652 -6027 -3628
rect -6013 -3658 -6012 -3634
rect -6010 -3658 -6008 -3634
rect -6004 -3658 -6002 -3634
rect -6000 -3658 -5999 -3634
rect -4289 -3651 -4288 -3611
rect -4286 -3651 -4285 -3611
rect -3799 -3647 -3798 -3635
rect -3796 -3647 -3795 -3635
rect -6080 -3691 -6079 -3679
rect -6077 -3691 -6076 -3679
rect -3760 -3663 -3759 -3639
rect -3757 -3663 -3755 -3639
rect -3751 -3663 -3749 -3639
rect -3747 -3663 -3746 -3639
rect -3732 -3669 -3731 -3645
rect -3729 -3669 -3727 -3645
rect -3723 -3669 -3721 -3645
rect -3719 -3669 -3718 -3645
rect -3799 -3702 -3798 -3690
rect -3796 -3702 -3795 -3690
rect -6077 -3780 -6076 -3768
rect -6074 -3780 -6073 -3768
rect -6038 -3796 -6037 -3772
rect -6035 -3796 -6033 -3772
rect -6029 -3796 -6027 -3772
rect -6025 -3796 -6024 -3772
rect -6010 -3802 -6009 -3778
rect -6007 -3802 -6005 -3778
rect -6001 -3802 -5999 -3778
rect -5997 -3802 -5996 -3778
rect -6077 -3835 -6076 -3823
rect -6074 -3835 -6073 -3823
rect -4290 -3794 -4289 -3754
rect -4287 -3794 -4286 -3754
rect -3798 -3790 -3797 -3778
rect -3795 -3790 -3794 -3778
rect -3759 -3806 -3758 -3782
rect -3756 -3806 -3754 -3782
rect -3750 -3806 -3748 -3782
rect -3746 -3806 -3745 -3782
rect -3731 -3812 -3730 -3788
rect -3728 -3812 -3726 -3788
rect -3722 -3812 -3720 -3788
rect -3718 -3812 -3717 -3788
rect -3798 -3845 -3797 -3833
rect -3795 -3845 -3794 -3833
rect -6081 -3928 -6080 -3916
rect -6078 -3928 -6077 -3916
rect -6042 -3944 -6041 -3920
rect -6039 -3944 -6037 -3920
rect -6033 -3944 -6031 -3920
rect -6029 -3944 -6028 -3920
rect -6014 -3950 -6013 -3926
rect -6011 -3950 -6009 -3926
rect -6005 -3950 -6003 -3926
rect -6001 -3950 -6000 -3926
rect -6081 -3983 -6080 -3971
rect -6078 -3983 -6077 -3971
rect -4290 -3946 -4289 -3906
rect -4287 -3946 -4286 -3906
rect -6056 -4144 -6055 -4132
rect -6053 -4144 -6052 -4132
rect -6017 -4160 -6016 -4136
rect -6014 -4160 -6012 -4136
rect -6008 -4160 -6006 -4136
rect -6004 -4160 -6003 -4136
rect -5989 -4166 -5988 -4142
rect -5986 -4166 -5984 -4142
rect -5980 -4166 -5978 -4142
rect -5976 -4166 -5975 -4142
rect -6056 -4199 -6055 -4187
rect -6053 -4199 -6052 -4187
rect -6057 -4395 -6056 -4375
rect -6054 -4395 -6050 -4375
rect -6046 -4395 -6045 -4375
rect -6043 -4395 -6042 -4375
rect -6015 -4402 -6014 -4382
rect -6012 -4402 -6011 -4382
rect -6056 -4504 -6055 -4484
rect -6053 -4504 -6049 -4484
rect -6045 -4504 -6044 -4484
rect -6042 -4504 -6041 -4484
rect -6014 -4511 -6013 -4491
rect -6011 -4511 -6010 -4491
rect -6053 -4632 -6052 -4612
rect -6050 -4632 -6046 -4612
rect -6042 -4632 -6041 -4612
rect -6039 -4632 -6038 -4612
rect -6011 -4639 -6010 -4619
rect -6008 -4639 -6007 -4619
rect -6051 -4752 -6050 -4732
rect -6048 -4752 -6044 -4732
rect -6040 -4752 -6039 -4732
rect -6037 -4752 -6036 -4732
rect -6009 -4759 -6008 -4739
rect -6006 -4759 -6005 -4739
rect -6049 -4893 -6048 -4873
rect -6046 -4893 -6042 -4873
rect -6038 -4893 -6037 -4873
rect -6035 -4893 -6034 -4873
rect -6007 -4900 -6006 -4880
rect -6004 -4900 -6003 -4880
rect -5227 -4912 -5226 -4872
rect -5224 -4912 -5223 -4872
<< ndcontact >>
rect -5237 -3068 -5233 -3048
rect -5229 -3068 -5225 -3048
rect -3733 -3225 -3729 -3219
rect -3725 -3225 -3721 -3219
rect -3694 -3274 -3690 -3262
rect -3676 -3274 -3672 -3262
rect -3666 -3274 -3662 -3262
rect -3648 -3274 -3644 -3262
rect -3733 -3280 -3729 -3274
rect -3725 -3280 -3721 -3274
rect -6077 -3484 -6073 -3478
rect -6069 -3484 -6065 -3478
rect -5095 -3499 -5091 -3399
rect -5087 -3499 -5083 -3399
rect -4294 -3427 -4290 -3407
rect -4286 -3427 -4282 -3407
rect -3802 -3409 -3798 -3403
rect -3794 -3409 -3790 -3403
rect -3763 -3458 -3759 -3446
rect -3745 -3458 -3741 -3446
rect -3735 -3458 -3731 -3446
rect -3717 -3458 -3713 -3446
rect -3802 -3464 -3798 -3458
rect -3794 -3464 -3790 -3458
rect -6038 -3533 -6034 -3521
rect -6020 -3533 -6016 -3521
rect -6010 -3533 -6006 -3521
rect -5992 -3533 -5988 -3521
rect -6077 -3539 -6073 -3533
rect -6069 -3539 -6065 -3533
rect -4923 -3588 -4919 -3488
rect -4915 -3588 -4911 -3488
rect -4293 -3558 -4289 -3538
rect -4285 -3558 -4281 -3538
rect -3807 -3539 -3803 -3533
rect -3799 -3539 -3795 -3533
rect -3768 -3588 -3764 -3576
rect -3750 -3588 -3746 -3576
rect -3740 -3588 -3736 -3576
rect -3722 -3588 -3718 -3576
rect -3807 -3594 -3803 -3588
rect -3799 -3594 -3795 -3588
rect -6084 -3656 -6080 -3650
rect -6076 -3656 -6072 -3650
rect -6045 -3705 -6041 -3693
rect -6027 -3705 -6023 -3693
rect -6017 -3705 -6013 -3693
rect -5999 -3705 -5995 -3693
rect -6084 -3711 -6080 -3705
rect -6076 -3711 -6072 -3705
rect -5087 -3767 -5083 -3667
rect -5079 -3767 -5075 -3667
rect -3803 -3667 -3799 -3661
rect -3795 -3667 -3791 -3661
rect -4293 -3689 -4289 -3669
rect -4285 -3689 -4281 -3669
rect -3764 -3716 -3760 -3704
rect -3746 -3716 -3742 -3704
rect -3736 -3716 -3732 -3704
rect -3718 -3716 -3714 -3704
rect -3803 -3722 -3799 -3716
rect -3795 -3722 -3791 -3716
rect -6081 -3800 -6077 -3794
rect -6073 -3800 -6069 -3794
rect -4749 -3822 -4745 -3722
rect -4741 -3822 -4737 -3722
rect -6042 -3849 -6038 -3837
rect -6024 -3849 -6020 -3837
rect -6014 -3849 -6010 -3837
rect -5996 -3849 -5992 -3837
rect -6081 -3855 -6077 -3849
rect -6073 -3855 -6069 -3849
rect -4625 -3853 -4621 -3753
rect -4617 -3853 -4613 -3753
rect -3802 -3810 -3798 -3804
rect -3794 -3810 -3790 -3804
rect -4294 -3832 -4290 -3812
rect -4286 -3832 -4282 -3812
rect -3763 -3859 -3759 -3847
rect -3745 -3859 -3741 -3847
rect -3735 -3859 -3731 -3847
rect -3717 -3859 -3713 -3847
rect -3802 -3865 -3798 -3859
rect -3794 -3865 -3790 -3859
rect -6085 -3948 -6081 -3942
rect -6077 -3948 -6073 -3942
rect -6046 -3997 -6042 -3985
rect -6028 -3997 -6024 -3985
rect -6018 -3997 -6014 -3985
rect -6000 -3997 -5996 -3985
rect -6085 -4003 -6081 -3997
rect -6077 -4003 -6073 -3997
rect -4485 -4016 -4481 -3916
rect -4477 -4016 -4473 -3916
rect -4294 -3984 -4290 -3964
rect -4286 -3984 -4282 -3964
rect -6060 -4164 -6056 -4158
rect -6052 -4164 -6048 -4158
rect -6021 -4213 -6017 -4201
rect -6003 -4213 -5999 -4201
rect -5993 -4213 -5989 -4201
rect -5975 -4213 -5971 -4201
rect -6060 -4219 -6056 -4213
rect -6052 -4219 -6048 -4213
rect -4914 -4391 -4910 -4291
rect -4906 -4391 -4902 -4291
rect -6061 -4444 -6057 -4424
rect -6042 -4444 -6038 -4424
rect -6019 -4426 -6015 -4416
rect -6011 -4426 -6007 -4416
rect -4740 -4424 -4736 -4324
rect -4732 -4424 -4728 -4324
rect -4616 -4495 -4612 -4395
rect -4608 -4495 -4604 -4395
rect -6060 -4553 -6056 -4533
rect -6041 -4553 -6037 -4533
rect -6018 -4535 -6014 -4525
rect -6010 -4535 -6006 -4525
rect -4477 -4594 -4473 -4494
rect -4469 -4594 -4465 -4494
rect -4398 -4653 -4394 -4553
rect -4390 -4653 -4386 -4553
rect -6057 -4681 -6053 -4661
rect -6038 -4681 -6034 -4661
rect -6015 -4663 -6011 -4653
rect -6007 -4663 -6003 -4653
rect -6055 -4801 -6051 -4781
rect -6036 -4801 -6032 -4781
rect -6013 -4783 -6009 -4773
rect -6005 -4783 -6001 -4773
rect -5078 -4911 -5074 -4811
rect -5070 -4911 -5066 -4811
rect -6053 -4942 -6049 -4922
rect -6034 -4942 -6030 -4922
rect -6011 -4924 -6007 -4914
rect -6003 -4924 -5999 -4914
rect -5231 -4950 -5227 -4930
rect -5223 -4950 -5219 -4930
<< pdcontact >>
rect -5237 -3030 -5233 -2990
rect -5229 -3030 -5225 -2990
rect -3733 -3205 -3729 -3193
rect -3725 -3205 -3721 -3193
rect -5103 -3267 -5099 -3217
rect -5095 -3267 -5091 -3217
rect -4931 -3268 -4927 -3218
rect -4923 -3268 -4919 -3218
rect -4757 -3268 -4753 -3218
rect -4749 -3268 -4745 -3218
rect -4633 -3269 -4629 -3219
rect -4625 -3269 -4621 -3219
rect -4493 -3272 -4489 -3222
rect -4485 -3272 -4481 -3222
rect -3694 -3221 -3690 -3197
rect -3685 -3221 -3681 -3197
rect -3676 -3221 -3672 -3197
rect -3666 -3227 -3662 -3203
rect -3657 -3227 -3653 -3203
rect -3648 -3227 -3644 -3203
rect -3733 -3260 -3729 -3248
rect -3725 -3260 -3721 -3248
rect -4294 -3389 -4290 -3349
rect -4286 -3389 -4282 -3349
rect -3802 -3389 -3798 -3377
rect -3794 -3389 -3790 -3377
rect -6077 -3464 -6073 -3452
rect -6069 -3464 -6065 -3452
rect -6038 -3480 -6034 -3456
rect -6029 -3480 -6025 -3456
rect -6020 -3480 -6016 -3456
rect -6010 -3486 -6006 -3462
rect -6001 -3486 -5997 -3462
rect -5992 -3486 -5988 -3462
rect -6077 -3519 -6073 -3507
rect -6069 -3519 -6065 -3507
rect -3763 -3405 -3759 -3381
rect -3754 -3405 -3750 -3381
rect -3745 -3405 -3741 -3381
rect -3735 -3411 -3731 -3387
rect -3726 -3411 -3722 -3387
rect -3717 -3411 -3713 -3387
rect -3802 -3444 -3798 -3432
rect -3794 -3444 -3790 -3432
rect -4293 -3520 -4289 -3480
rect -4285 -3520 -4281 -3480
rect -3807 -3519 -3803 -3507
rect -3799 -3519 -3795 -3507
rect -3768 -3535 -3764 -3511
rect -3759 -3535 -3755 -3511
rect -3750 -3535 -3746 -3511
rect -3740 -3541 -3736 -3517
rect -3731 -3541 -3727 -3517
rect -3722 -3541 -3718 -3517
rect -3807 -3574 -3803 -3562
rect -3799 -3574 -3795 -3562
rect -6084 -3636 -6080 -3624
rect -6076 -3636 -6072 -3624
rect -6045 -3652 -6041 -3628
rect -6036 -3652 -6032 -3628
rect -6027 -3652 -6023 -3628
rect -6017 -3658 -6013 -3634
rect -6008 -3658 -6004 -3634
rect -5999 -3658 -5995 -3634
rect -4293 -3651 -4289 -3611
rect -4285 -3651 -4281 -3611
rect -3803 -3647 -3799 -3635
rect -3795 -3647 -3791 -3635
rect -6084 -3691 -6080 -3679
rect -6076 -3691 -6072 -3679
rect -3764 -3663 -3760 -3639
rect -3755 -3663 -3751 -3639
rect -3746 -3663 -3742 -3639
rect -3736 -3669 -3732 -3645
rect -3727 -3669 -3723 -3645
rect -3718 -3669 -3714 -3645
rect -3803 -3702 -3799 -3690
rect -3795 -3702 -3791 -3690
rect -6081 -3780 -6077 -3768
rect -6073 -3780 -6069 -3768
rect -6042 -3796 -6038 -3772
rect -6033 -3796 -6029 -3772
rect -6024 -3796 -6020 -3772
rect -6014 -3802 -6010 -3778
rect -6005 -3802 -6001 -3778
rect -5996 -3802 -5992 -3778
rect -6081 -3835 -6077 -3823
rect -6073 -3835 -6069 -3823
rect -4294 -3794 -4290 -3754
rect -4286 -3794 -4282 -3754
rect -3802 -3790 -3798 -3778
rect -3794 -3790 -3790 -3778
rect -3763 -3806 -3759 -3782
rect -3754 -3806 -3750 -3782
rect -3745 -3806 -3741 -3782
rect -3735 -3812 -3731 -3788
rect -3726 -3812 -3722 -3788
rect -3717 -3812 -3713 -3788
rect -3802 -3845 -3798 -3833
rect -3794 -3845 -3790 -3833
rect -6085 -3928 -6081 -3916
rect -6077 -3928 -6073 -3916
rect -6046 -3944 -6042 -3920
rect -6037 -3944 -6033 -3920
rect -6028 -3944 -6024 -3920
rect -6018 -3950 -6014 -3926
rect -6009 -3950 -6005 -3926
rect -6000 -3950 -5996 -3926
rect -6085 -3983 -6081 -3971
rect -6077 -3983 -6073 -3971
rect -4294 -3946 -4290 -3906
rect -4286 -3946 -4282 -3906
rect -6060 -4144 -6056 -4132
rect -6052 -4144 -6048 -4132
rect -6021 -4160 -6017 -4136
rect -6012 -4160 -6008 -4136
rect -6003 -4160 -5999 -4136
rect -5993 -4166 -5989 -4142
rect -5984 -4166 -5980 -4142
rect -5975 -4166 -5971 -4142
rect -6060 -4199 -6056 -4187
rect -6052 -4199 -6048 -4187
rect -6061 -4395 -6057 -4375
rect -6050 -4395 -6046 -4375
rect -6042 -4395 -6038 -4375
rect -6019 -4402 -6015 -4382
rect -6011 -4402 -6007 -4382
rect -6060 -4504 -6056 -4484
rect -6049 -4504 -6045 -4484
rect -6041 -4504 -6037 -4484
rect -6018 -4511 -6014 -4491
rect -6010 -4511 -6006 -4491
rect -6057 -4632 -6053 -4612
rect -6046 -4632 -6042 -4612
rect -6038 -4632 -6034 -4612
rect -6015 -4639 -6011 -4619
rect -6007 -4639 -6003 -4619
rect -6055 -4752 -6051 -4732
rect -6044 -4752 -6040 -4732
rect -6036 -4752 -6032 -4732
rect -6013 -4759 -6009 -4739
rect -6005 -4759 -6001 -4739
rect -6053 -4893 -6049 -4873
rect -6042 -4893 -6038 -4873
rect -6034 -4893 -6030 -4873
rect -6011 -4900 -6007 -4880
rect -6003 -4900 -5999 -4880
rect -5231 -4912 -5227 -4872
rect -5223 -4912 -5219 -4872
<< psubstratepcontact >>
rect -6005 -4435 -6000 -4431
rect -6004 -4544 -5999 -4540
rect -6001 -4672 -5996 -4668
rect -5999 -4792 -5994 -4788
rect -5997 -4933 -5992 -4929
<< nsubstratencontact >>
rect -5242 -2984 -5238 -2980
rect -5108 -3211 -5104 -3206
rect -4936 -3212 -4932 -3207
rect -4762 -3212 -4758 -3207
rect -4638 -3213 -4634 -3208
rect -4498 -3216 -4494 -3211
rect -4299 -3343 -4295 -3339
rect -4298 -3474 -4294 -3470
rect -4298 -3605 -4294 -3601
rect -4299 -3748 -4295 -3744
rect -4299 -3900 -4295 -3896
rect -6061 -4370 -6057 -4364
rect -6009 -4375 -6005 -4371
rect -6060 -4479 -6056 -4473
rect -6008 -4484 -6004 -4480
rect -6057 -4607 -6053 -4601
rect -6005 -4612 -6001 -4608
rect -6055 -4727 -6051 -4721
rect -6003 -4732 -5999 -4728
rect -6053 -4868 -6049 -4862
rect -5236 -4866 -5232 -4862
rect -6001 -4873 -5997 -4869
<< polysilicon >>
rect -5232 -2990 -5230 -2987
rect -5232 -3048 -5230 -3030
rect -5232 -3072 -5230 -3068
rect -3728 -3193 -3726 -3190
rect -3689 -3197 -3687 -3194
rect -3679 -3197 -3677 -3194
rect -5098 -3217 -5096 -3214
rect -4926 -3218 -4924 -3215
rect -4752 -3218 -4750 -3215
rect -5098 -3290 -5096 -3267
rect -4628 -3219 -4626 -3216
rect -3728 -3219 -3726 -3205
rect -4926 -3291 -4924 -3268
rect -4752 -3291 -4750 -3268
rect -4488 -3222 -4486 -3219
rect -4628 -3292 -4626 -3269
rect -3661 -3203 -3659 -3200
rect -3651 -3203 -3649 -3200
rect -3728 -3228 -3726 -3225
rect -3689 -3230 -3687 -3221
rect -3679 -3231 -3677 -3221
rect -3728 -3248 -3726 -3245
rect -4488 -3295 -4486 -3272
rect -3728 -3274 -3726 -3260
rect -3689 -3262 -3687 -3235
rect -3679 -3262 -3677 -3236
rect -3661 -3238 -3659 -3227
rect -3661 -3262 -3659 -3242
rect -3651 -3249 -3649 -3227
rect -3651 -3262 -3649 -3253
rect -3689 -3277 -3687 -3274
rect -3679 -3277 -3677 -3274
rect -3661 -3277 -3659 -3274
rect -3651 -3277 -3649 -3274
rect -3728 -3283 -3726 -3280
rect -4289 -3349 -4287 -3346
rect -3797 -3377 -3795 -3374
rect -3758 -3381 -3756 -3378
rect -3748 -3381 -3746 -3378
rect -5090 -3399 -5088 -3396
rect -6072 -3452 -6070 -3449
rect -6033 -3456 -6031 -3453
rect -6023 -3456 -6021 -3453
rect -6072 -3478 -6070 -3464
rect -6005 -3462 -6003 -3459
rect -5995 -3462 -5993 -3459
rect -6072 -3487 -6070 -3484
rect -6033 -3489 -6031 -3480
rect -6023 -3490 -6021 -3480
rect -6072 -3507 -6070 -3504
rect -6072 -3533 -6070 -3519
rect -6033 -3521 -6031 -3494
rect -6023 -3521 -6021 -3495
rect -6005 -3497 -6003 -3486
rect -6005 -3521 -6003 -3501
rect -5995 -3508 -5993 -3486
rect -4289 -3407 -4287 -3389
rect -3797 -3403 -3795 -3389
rect -3730 -3387 -3728 -3384
rect -3720 -3387 -3718 -3384
rect -3797 -3412 -3795 -3409
rect -3758 -3414 -3756 -3405
rect -3748 -3415 -3746 -3405
rect -4289 -3431 -4287 -3427
rect -3797 -3432 -3795 -3429
rect -3797 -3458 -3795 -3444
rect -3758 -3446 -3756 -3419
rect -3748 -3446 -3746 -3420
rect -3730 -3422 -3728 -3411
rect -3730 -3446 -3728 -3426
rect -3720 -3433 -3718 -3411
rect -3720 -3446 -3718 -3437
rect -3758 -3461 -3756 -3458
rect -3748 -3461 -3746 -3458
rect -3730 -3461 -3728 -3458
rect -3720 -3461 -3718 -3458
rect -3797 -3467 -3795 -3464
rect -4288 -3480 -4286 -3477
rect -4918 -3488 -4916 -3485
rect -5995 -3521 -5993 -3512
rect -5090 -3515 -5088 -3499
rect -6033 -3536 -6031 -3533
rect -6023 -3536 -6021 -3533
rect -6005 -3536 -6003 -3533
rect -5995 -3536 -5993 -3533
rect -6072 -3542 -6070 -3539
rect -3802 -3507 -3800 -3504
rect -3763 -3511 -3761 -3508
rect -3753 -3511 -3751 -3508
rect -4288 -3538 -4286 -3520
rect -3802 -3533 -3800 -3519
rect -3735 -3517 -3733 -3514
rect -3725 -3517 -3723 -3514
rect -3802 -3542 -3800 -3539
rect -3763 -3544 -3761 -3535
rect -3753 -3545 -3751 -3535
rect -4288 -3562 -4286 -3558
rect -3802 -3562 -3800 -3559
rect -3802 -3588 -3800 -3574
rect -3763 -3576 -3761 -3549
rect -3753 -3576 -3751 -3550
rect -3735 -3552 -3733 -3541
rect -3735 -3576 -3733 -3556
rect -3725 -3563 -3723 -3541
rect -3725 -3576 -3723 -3567
rect -4918 -3604 -4916 -3588
rect -3763 -3591 -3761 -3588
rect -3753 -3591 -3751 -3588
rect -3735 -3591 -3733 -3588
rect -3725 -3591 -3723 -3588
rect -3802 -3597 -3800 -3594
rect -4288 -3611 -4286 -3608
rect -6079 -3624 -6077 -3621
rect -6040 -3628 -6038 -3625
rect -6030 -3628 -6028 -3625
rect -6079 -3650 -6077 -3636
rect -6012 -3634 -6010 -3631
rect -6002 -3634 -6000 -3631
rect -6079 -3659 -6077 -3656
rect -6040 -3661 -6038 -3652
rect -6030 -3662 -6028 -3652
rect -3798 -3635 -3796 -3632
rect -3759 -3639 -3757 -3636
rect -3749 -3639 -3747 -3636
rect -6079 -3679 -6077 -3676
rect -6079 -3705 -6077 -3691
rect -6040 -3693 -6038 -3666
rect -6030 -3693 -6028 -3667
rect -6012 -3669 -6010 -3658
rect -6012 -3693 -6010 -3673
rect -6002 -3680 -6000 -3658
rect -5082 -3667 -5080 -3664
rect -6002 -3693 -6000 -3684
rect -6040 -3708 -6038 -3705
rect -6030 -3708 -6028 -3705
rect -6012 -3708 -6010 -3705
rect -6002 -3708 -6000 -3705
rect -6079 -3714 -6077 -3711
rect -6076 -3768 -6074 -3765
rect -4288 -3669 -4286 -3651
rect -3798 -3661 -3796 -3647
rect -3731 -3645 -3729 -3642
rect -3721 -3645 -3719 -3642
rect -3798 -3670 -3796 -3667
rect -3759 -3672 -3757 -3663
rect -3749 -3673 -3747 -3663
rect -4288 -3693 -4286 -3689
rect -3798 -3690 -3796 -3687
rect -3798 -3716 -3796 -3702
rect -3759 -3704 -3757 -3677
rect -3749 -3704 -3747 -3678
rect -3731 -3680 -3729 -3669
rect -3731 -3704 -3729 -3684
rect -3721 -3691 -3719 -3669
rect -3721 -3704 -3719 -3695
rect -4744 -3722 -4742 -3719
rect -3759 -3719 -3757 -3716
rect -3749 -3719 -3747 -3716
rect -3731 -3719 -3729 -3716
rect -3721 -3719 -3719 -3716
rect -6037 -3772 -6035 -3769
rect -6027 -3772 -6025 -3769
rect -6076 -3794 -6074 -3780
rect -6009 -3778 -6007 -3775
rect -5999 -3778 -5997 -3775
rect -6076 -3803 -6074 -3800
rect -6037 -3805 -6035 -3796
rect -6027 -3806 -6025 -3796
rect -5082 -3783 -5080 -3767
rect -6076 -3823 -6074 -3820
rect -6076 -3849 -6074 -3835
rect -6037 -3837 -6035 -3810
rect -6027 -3837 -6025 -3811
rect -6009 -3813 -6007 -3802
rect -6009 -3837 -6007 -3817
rect -5999 -3824 -5997 -3802
rect -3798 -3725 -3796 -3722
rect -4620 -3753 -4618 -3750
rect -5999 -3837 -5997 -3828
rect -4744 -3838 -4742 -3822
rect -6037 -3852 -6035 -3849
rect -6027 -3852 -6025 -3849
rect -6009 -3852 -6007 -3849
rect -5999 -3852 -5997 -3849
rect -4289 -3754 -4287 -3751
rect -3797 -3778 -3795 -3775
rect -3758 -3782 -3756 -3779
rect -3748 -3782 -3746 -3779
rect -4289 -3812 -4287 -3794
rect -3797 -3804 -3795 -3790
rect -3730 -3788 -3728 -3785
rect -3720 -3788 -3718 -3785
rect -3797 -3813 -3795 -3810
rect -3758 -3815 -3756 -3806
rect -3748 -3816 -3746 -3806
rect -4289 -3836 -4287 -3832
rect -3797 -3833 -3795 -3830
rect -6076 -3858 -6074 -3855
rect -4620 -3869 -4618 -3853
rect -3797 -3859 -3795 -3845
rect -3758 -3847 -3756 -3820
rect -3748 -3847 -3746 -3821
rect -3730 -3823 -3728 -3812
rect -3730 -3847 -3728 -3827
rect -3720 -3834 -3718 -3812
rect -3720 -3847 -3718 -3838
rect -3758 -3862 -3756 -3859
rect -3748 -3862 -3746 -3859
rect -3730 -3862 -3728 -3859
rect -3720 -3862 -3718 -3859
rect -3797 -3868 -3795 -3865
rect -4289 -3906 -4287 -3903
rect -6080 -3916 -6078 -3913
rect -4480 -3916 -4478 -3913
rect -6041 -3920 -6039 -3917
rect -6031 -3920 -6029 -3917
rect -6080 -3942 -6078 -3928
rect -6013 -3926 -6011 -3923
rect -6003 -3926 -6001 -3923
rect -6080 -3951 -6078 -3948
rect -6041 -3953 -6039 -3944
rect -6031 -3954 -6029 -3944
rect -6080 -3971 -6078 -3968
rect -6080 -3997 -6078 -3983
rect -6041 -3985 -6039 -3958
rect -6031 -3985 -6029 -3959
rect -6013 -3961 -6011 -3950
rect -6013 -3985 -6011 -3965
rect -6003 -3972 -6001 -3950
rect -6003 -3985 -6001 -3976
rect -6041 -4000 -6039 -3997
rect -6031 -4000 -6029 -3997
rect -6013 -4000 -6011 -3997
rect -6003 -4000 -6001 -3997
rect -6080 -4006 -6078 -4003
rect -4289 -3964 -4287 -3946
rect -4289 -3988 -4287 -3984
rect -4480 -4032 -4478 -4016
rect -6055 -4132 -6053 -4129
rect -6016 -4136 -6014 -4133
rect -6006 -4136 -6004 -4133
rect -6055 -4158 -6053 -4144
rect -5988 -4142 -5986 -4139
rect -5978 -4142 -5976 -4139
rect -6055 -4167 -6053 -4164
rect -6016 -4169 -6014 -4160
rect -6006 -4170 -6004 -4160
rect -6055 -4187 -6053 -4184
rect -6055 -4213 -6053 -4199
rect -6016 -4201 -6014 -4174
rect -6006 -4201 -6004 -4175
rect -5988 -4177 -5986 -4166
rect -5988 -4201 -5986 -4181
rect -5978 -4188 -5976 -4166
rect -5978 -4201 -5976 -4192
rect -6016 -4216 -6014 -4213
rect -6006 -4216 -6004 -4213
rect -5988 -4216 -5986 -4213
rect -5978 -4216 -5976 -4213
rect -6055 -4222 -6053 -4219
rect -4909 -4291 -4907 -4288
rect -6056 -4375 -6054 -4372
rect -6045 -4375 -6043 -4372
rect -6014 -4382 -6012 -4378
rect -6056 -4424 -6054 -4395
rect -6045 -4424 -6043 -4395
rect -4735 -4324 -4733 -4321
rect -6014 -4416 -6012 -4402
rect -4909 -4407 -4907 -4391
rect -4611 -4395 -4609 -4392
rect -6014 -4429 -6012 -4426
rect -4735 -4440 -4733 -4424
rect -6056 -4447 -6054 -4444
rect -6045 -4447 -6043 -4444
rect -6055 -4484 -6053 -4481
rect -6044 -4484 -6042 -4481
rect -6013 -4491 -6011 -4487
rect -6055 -4533 -6053 -4504
rect -6044 -4533 -6042 -4504
rect -4472 -4494 -4470 -4491
rect -4611 -4511 -4609 -4495
rect -6013 -4525 -6011 -4511
rect -6013 -4538 -6011 -4535
rect -6055 -4556 -6053 -4553
rect -6044 -4556 -6042 -4553
rect -4393 -4553 -4391 -4550
rect -6052 -4612 -6050 -4609
rect -6041 -4612 -6039 -4609
rect -4472 -4610 -4470 -4594
rect -6010 -4619 -6008 -4615
rect -6052 -4661 -6050 -4632
rect -6041 -4661 -6039 -4632
rect -6010 -4653 -6008 -4639
rect -6010 -4666 -6008 -4663
rect -4393 -4669 -4391 -4653
rect -6052 -4684 -6050 -4681
rect -6041 -4684 -6039 -4681
rect -6050 -4732 -6048 -4729
rect -6039 -4732 -6037 -4729
rect -6008 -4739 -6006 -4735
rect -6050 -4781 -6048 -4752
rect -6039 -4781 -6037 -4752
rect -6008 -4773 -6006 -4759
rect -6008 -4786 -6006 -4783
rect -6050 -4804 -6048 -4801
rect -6039 -4804 -6037 -4801
rect -5073 -4811 -5071 -4808
rect -6048 -4873 -6046 -4870
rect -6037 -4873 -6035 -4870
rect -5226 -4872 -5224 -4869
rect -6006 -4880 -6004 -4876
rect -6048 -4922 -6046 -4893
rect -6037 -4922 -6035 -4893
rect -6006 -4914 -6004 -4900
rect -6006 -4927 -6004 -4924
rect -5226 -4930 -5224 -4912
rect -5073 -4927 -5071 -4911
rect -6048 -4945 -6046 -4942
rect -6037 -4945 -6035 -4942
rect -5226 -4954 -5224 -4950
<< polycontact >>
rect -3732 -3216 -3728 -3212
rect -3732 -3271 -3728 -3267
rect -3663 -3242 -3659 -3238
rect -3652 -3253 -3648 -3249
rect -6076 -3475 -6072 -3471
rect -6076 -3530 -6072 -3526
rect -6007 -3501 -6003 -3497
rect -3801 -3400 -3797 -3396
rect -3801 -3455 -3797 -3451
rect -3732 -3426 -3728 -3422
rect -3721 -3437 -3717 -3433
rect -5996 -3512 -5992 -3508
rect -3806 -3530 -3802 -3526
rect -3806 -3585 -3802 -3581
rect -3737 -3556 -3733 -3552
rect -3726 -3567 -3722 -3563
rect -6083 -3647 -6079 -3643
rect -6083 -3702 -6079 -3698
rect -6014 -3673 -6010 -3669
rect -6003 -3684 -5999 -3680
rect -3802 -3658 -3798 -3654
rect -3802 -3713 -3798 -3709
rect -3733 -3684 -3729 -3680
rect -3722 -3695 -3718 -3691
rect -6080 -3791 -6076 -3787
rect -6080 -3846 -6076 -3842
rect -6011 -3817 -6007 -3813
rect -6000 -3828 -5996 -3824
rect -3801 -3801 -3797 -3797
rect -3801 -3856 -3797 -3852
rect -3732 -3827 -3728 -3823
rect -3721 -3838 -3717 -3834
rect -6084 -3939 -6080 -3935
rect -6084 -3994 -6080 -3990
rect -6015 -3965 -6011 -3961
rect -6004 -3976 -6000 -3972
rect -6059 -4155 -6055 -4151
rect -6059 -4210 -6055 -4206
rect -5990 -4181 -5986 -4177
rect -5979 -4192 -5975 -4188
rect -6060 -4421 -6056 -4417
rect -6049 -4414 -6045 -4410
rect -6018 -4413 -6014 -4409
rect -6059 -4530 -6055 -4526
rect -6048 -4523 -6044 -4519
rect -6017 -4522 -6013 -4518
rect -6056 -4658 -6052 -4654
rect -6045 -4651 -6041 -4647
rect -6014 -4650 -6010 -4646
rect -6054 -4778 -6050 -4774
rect -6043 -4771 -6039 -4767
rect -6012 -4770 -6008 -4766
rect -6052 -4919 -6048 -4915
rect -6041 -4912 -6037 -4908
rect -6010 -4911 -6006 -4907
<< metal1 >>
rect -5882 -3169 -5877 -2602
rect -6316 -3174 -5877 -3169
rect -6078 -3446 -6050 -3443
rect -6077 -3452 -6074 -3446
rect -6053 -3447 -6050 -3446
rect -6053 -3450 -5982 -3447
rect -6288 -3476 -6091 -3473
rect -6086 -3475 -6076 -3472
rect -6068 -3472 -6065 -3464
rect -6038 -3456 -6035 -3450
rect -6019 -3456 -6016 -3450
rect -6068 -3475 -6047 -3472
rect -6068 -3478 -6065 -3475
rect -6077 -3488 -6074 -3484
rect -6083 -3490 -6059 -3488
rect -6083 -3491 -6065 -3490
rect -6060 -3491 -6059 -3490
rect -6050 -3498 -6047 -3475
rect -6009 -3456 -5989 -3453
rect -6009 -3462 -6006 -3456
rect -5992 -3462 -5989 -3456
rect -6028 -3483 -6025 -3480
rect -6028 -3486 -6010 -3483
rect -6000 -3493 -5997 -3486
rect -6000 -3496 -5983 -3493
rect -6078 -3499 -6059 -3498
rect -6083 -3501 -6059 -3499
rect -6050 -3501 -6007 -3498
rect -6077 -3507 -6074 -3501
rect -5986 -3507 -5983 -3496
rect -6021 -3512 -5996 -3509
rect -5986 -3510 -5972 -3507
rect -5986 -3511 -5977 -3510
rect -6021 -3514 -6018 -3512
rect -6271 -3530 -6091 -3527
rect -6086 -3530 -6076 -3527
rect -6068 -3527 -6065 -3519
rect -6056 -3517 -6018 -3514
rect -5986 -3515 -5983 -3511
rect -6056 -3527 -6053 -3517
rect -6015 -3518 -5983 -3515
rect -6015 -3521 -6012 -3518
rect -6068 -3530 -6053 -3527
rect -6068 -3533 -6065 -3530
rect -6016 -3524 -6010 -3521
rect -6077 -3543 -6074 -3539
rect -6056 -3540 -6051 -3537
rect -6038 -3537 -6035 -3533
rect -5991 -3537 -5988 -3533
rect -6046 -3540 -5982 -3537
rect -6056 -3543 -6053 -3540
rect -6083 -3546 -6053 -3543
rect -6085 -3618 -6057 -3615
rect -6084 -3624 -6081 -3618
rect -6060 -3619 -6057 -3618
rect -6060 -3622 -5989 -3619
rect -6181 -3648 -6098 -3645
rect -6093 -3647 -6083 -3644
rect -6075 -3644 -6072 -3636
rect -6045 -3628 -6042 -3622
rect -6026 -3628 -6023 -3622
rect -6075 -3647 -6054 -3644
rect -6075 -3650 -6072 -3647
rect -6084 -3660 -6081 -3656
rect -6090 -3662 -6066 -3660
rect -6090 -3663 -6072 -3662
rect -6067 -3663 -6066 -3662
rect -6057 -3670 -6054 -3647
rect -6016 -3628 -5996 -3625
rect -6016 -3634 -6013 -3628
rect -5999 -3634 -5996 -3628
rect -6035 -3655 -6032 -3652
rect -6035 -3658 -6017 -3655
rect -6007 -3665 -6004 -3658
rect -6007 -3668 -5990 -3665
rect -6085 -3671 -6066 -3670
rect -6090 -3673 -6066 -3671
rect -6057 -3673 -6014 -3670
rect -6084 -3679 -6081 -3673
rect -5993 -3679 -5990 -3668
rect -5984 -3679 -5979 -3604
rect -6028 -3684 -6003 -3681
rect -5993 -3683 -5979 -3679
rect -6028 -3686 -6025 -3684
rect -6180 -3702 -6098 -3699
rect -6093 -3702 -6083 -3699
rect -6075 -3699 -6072 -3691
rect -6063 -3689 -6025 -3686
rect -5993 -3687 -5990 -3683
rect -6063 -3699 -6060 -3689
rect -6022 -3690 -5990 -3687
rect -6022 -3693 -6019 -3690
rect -6075 -3702 -6060 -3699
rect -6075 -3705 -6072 -3702
rect -6023 -3696 -6017 -3693
rect -6084 -3715 -6081 -3711
rect -6063 -3712 -6058 -3709
rect -6045 -3709 -6042 -3705
rect -5998 -3709 -5995 -3705
rect -6053 -3712 -5989 -3709
rect -6063 -3715 -6060 -3712
rect -6090 -3718 -6060 -3715
rect -6082 -3762 -6054 -3759
rect -6081 -3768 -6078 -3762
rect -6057 -3763 -6054 -3762
rect -6057 -3766 -5986 -3763
rect -6171 -3792 -6095 -3789
rect -6090 -3791 -6080 -3788
rect -6072 -3788 -6069 -3780
rect -6042 -3772 -6039 -3766
rect -6023 -3772 -6020 -3766
rect -6072 -3791 -6051 -3788
rect -6072 -3794 -6069 -3791
rect -6081 -3804 -6078 -3800
rect -6087 -3806 -6063 -3804
rect -6087 -3807 -6069 -3806
rect -6064 -3807 -6063 -3806
rect -6054 -3814 -6051 -3791
rect -6013 -3772 -5993 -3769
rect -6013 -3778 -6010 -3772
rect -5996 -3778 -5993 -3772
rect -5882 -3778 -5877 -3174
rect -5765 -3510 -5760 -2666
rect -5708 -3599 -5703 -2752
rect -6032 -3799 -6029 -3796
rect -6032 -3802 -6014 -3799
rect -6004 -3809 -6001 -3802
rect -6004 -3812 -5987 -3809
rect -6082 -3815 -6063 -3814
rect -6087 -3817 -6063 -3815
rect -6054 -3817 -6011 -3814
rect -6081 -3823 -6078 -3817
rect -5990 -3823 -5987 -3812
rect -6025 -3828 -6000 -3825
rect -5990 -3827 -5976 -3823
rect -6025 -3830 -6022 -3828
rect -6178 -3846 -6095 -3843
rect -6090 -3846 -6080 -3843
rect -6072 -3843 -6069 -3835
rect -6060 -3833 -6022 -3830
rect -5990 -3831 -5987 -3827
rect -6060 -3843 -6057 -3833
rect -6019 -3834 -5987 -3831
rect -5981 -3833 -5976 -3827
rect -6019 -3837 -6016 -3834
rect -6072 -3846 -6057 -3843
rect -6072 -3849 -6069 -3846
rect -6020 -3840 -6014 -3837
rect -5616 -3833 -5611 -2813
rect -6081 -3859 -6078 -3855
rect -6060 -3856 -6055 -3853
rect -6042 -3853 -6039 -3849
rect -5995 -3853 -5992 -3849
rect -6050 -3856 -5986 -3853
rect -6060 -3859 -6057 -3856
rect -6087 -3862 -6057 -3859
rect -5487 -3864 -5482 -2902
rect -6086 -3910 -6058 -3907
rect -6085 -3916 -6082 -3910
rect -6061 -3911 -6058 -3910
rect -6061 -3914 -5990 -3911
rect -6174 -3940 -6099 -3937
rect -6094 -3939 -6084 -3936
rect -6076 -3936 -6073 -3928
rect -6046 -3920 -6043 -3914
rect -6027 -3920 -6024 -3914
rect -6076 -3939 -6055 -3936
rect -6076 -3942 -6073 -3939
rect -6085 -3952 -6082 -3948
rect -6091 -3954 -6067 -3952
rect -6091 -3955 -6073 -3954
rect -6068 -3955 -6067 -3954
rect -6058 -3962 -6055 -3939
rect -6017 -3920 -5997 -3917
rect -6017 -3926 -6014 -3920
rect -6000 -3926 -5997 -3920
rect -6036 -3947 -6033 -3944
rect -6036 -3950 -6018 -3947
rect -6008 -3957 -6005 -3950
rect -6008 -3960 -5991 -3957
rect -6086 -3963 -6067 -3962
rect -6091 -3965 -6067 -3963
rect -6058 -3965 -6015 -3962
rect -6085 -3971 -6082 -3965
rect -5994 -3971 -5991 -3960
rect -5985 -3971 -5980 -3869
rect -6029 -3976 -6004 -3973
rect -5994 -3975 -5980 -3971
rect -6029 -3978 -6026 -3976
rect -6174 -3994 -6099 -3991
rect -6094 -3994 -6084 -3991
rect -6076 -3991 -6073 -3983
rect -6064 -3981 -6026 -3978
rect -5994 -3979 -5991 -3975
rect -6064 -3991 -6061 -3981
rect -6023 -3982 -5991 -3979
rect -6023 -3985 -6020 -3982
rect -6076 -3994 -6061 -3991
rect -6076 -3997 -6073 -3994
rect -6024 -3988 -6018 -3985
rect -6085 -4007 -6082 -4003
rect -6064 -4004 -6059 -4001
rect -6046 -4001 -6043 -3997
rect -5999 -4001 -5996 -3997
rect -6054 -4004 -5990 -4001
rect -6064 -4007 -6061 -4004
rect -6091 -4010 -6061 -4007
rect -5327 -4027 -5322 -2947
rect -5237 -2980 -5233 -2977
rect -5243 -2984 -5242 -2980
rect -5238 -2984 -5233 -2980
rect -5237 -2990 -5233 -2984
rect -5229 -3040 -5225 -3030
rect -5229 -3046 -5189 -3040
rect -5229 -3048 -5225 -3046
rect -5237 -3078 -5233 -3068
rect -5196 -3151 -5189 -3046
rect -5196 -3154 -4684 -3151
rect -5196 -3157 -4544 -3154
rect -5196 -3284 -5189 -3157
rect -5103 -3206 -5099 -3197
rect -5109 -3211 -5108 -3206
rect -5104 -3211 -5085 -3206
rect -5103 -3217 -5099 -3211
rect -5196 -3290 -5115 -3284
rect -5196 -3292 -5189 -3290
rect -5095 -3320 -5091 -3267
rect -4981 -3285 -4974 -3157
rect -4931 -3207 -4927 -3198
rect -4937 -3212 -4936 -3207
rect -4932 -3212 -4913 -3207
rect -4931 -3218 -4927 -3212
rect -4981 -3291 -4942 -3285
rect -5095 -3325 -4992 -3320
rect -5095 -3399 -5091 -3325
rect -4997 -3399 -4992 -3325
rect -5087 -3667 -5083 -3499
rect -4997 -3637 -4992 -3404
rect -4923 -3327 -4919 -3268
rect -4811 -3285 -4805 -3157
rect -4690 -3160 -4544 -3157
rect -4757 -3207 -4753 -3198
rect -4763 -3212 -4762 -3207
rect -4758 -3212 -4739 -3207
rect -4757 -3218 -4753 -3212
rect -4811 -3291 -4768 -3285
rect -4749 -3322 -4745 -3268
rect -4690 -3286 -4684 -3160
rect -4633 -3208 -4629 -3199
rect -4639 -3213 -4638 -3208
rect -4634 -3213 -4615 -3208
rect -4633 -3219 -4629 -3213
rect -4690 -3292 -4644 -3286
rect -4749 -3327 -4652 -3322
rect -4923 -3332 -4809 -3327
rect -4923 -3488 -4919 -3332
rect -4915 -3637 -4911 -3588
rect -4997 -3644 -4911 -3637
rect -6061 -4126 -6033 -4123
rect -6060 -4132 -6057 -4126
rect -6036 -4127 -6033 -4126
rect -6036 -4130 -5965 -4127
rect -6149 -4156 -6074 -4153
rect -6069 -4155 -6059 -4152
rect -6051 -4152 -6048 -4144
rect -6021 -4136 -6018 -4130
rect -6002 -4136 -5999 -4130
rect -6051 -4155 -6030 -4152
rect -6051 -4158 -6048 -4155
rect -6060 -4168 -6057 -4164
rect -6066 -4170 -6042 -4168
rect -6066 -4171 -6048 -4170
rect -6043 -4171 -6042 -4170
rect -6033 -4178 -6030 -4155
rect -5992 -4136 -5972 -4133
rect -5992 -4142 -5989 -4136
rect -5975 -4142 -5972 -4136
rect -6011 -4163 -6008 -4160
rect -6011 -4166 -5993 -4163
rect -5983 -4173 -5980 -4166
rect -5983 -4176 -5966 -4173
rect -6061 -4179 -6042 -4178
rect -6066 -4181 -6042 -4179
rect -6033 -4181 -5990 -4178
rect -6060 -4187 -6057 -4181
rect -5969 -4187 -5966 -4176
rect -5960 -4187 -5955 -4032
rect -6004 -4192 -5979 -4189
rect -5969 -4191 -5955 -4187
rect -6004 -4194 -6001 -4192
rect -6149 -4210 -6074 -4207
rect -6069 -4210 -6059 -4207
rect -6051 -4207 -6048 -4199
rect -6039 -4197 -6001 -4194
rect -5969 -4195 -5966 -4191
rect -6039 -4207 -6036 -4197
rect -5998 -4198 -5966 -4195
rect -5998 -4201 -5995 -4198
rect -6051 -4210 -6036 -4207
rect -6051 -4213 -6048 -4210
rect -5999 -4204 -5993 -4201
rect -6060 -4223 -6057 -4219
rect -6039 -4220 -6034 -4217
rect -6021 -4217 -6018 -4213
rect -5974 -4217 -5971 -4213
rect -6029 -4220 -5965 -4217
rect -6039 -4223 -6036 -4220
rect -6066 -4226 -6036 -4223
rect -5079 -4269 -5075 -3767
rect -4915 -4269 -4911 -3644
rect -4814 -3530 -4809 -3332
rect -4814 -3891 -4809 -3535
rect -4749 -3722 -4745 -3327
rect -4657 -3661 -4652 -3327
rect -4741 -3891 -4737 -3822
rect -4814 -3896 -4737 -3891
rect -4741 -4269 -4737 -3896
rect -4657 -3903 -4652 -3666
rect -4625 -3359 -4621 -3269
rect -4550 -3289 -4544 -3160
rect -4493 -3211 -4489 -3202
rect -4499 -3216 -4498 -3211
rect -4494 -3216 -4475 -3211
rect -4493 -3222 -4489 -3216
rect -4550 -3295 -4504 -3289
rect -4485 -3359 -4481 -3272
rect -4294 -3339 -4290 -3336
rect -4300 -3343 -4299 -3339
rect -4295 -3343 -4290 -3339
rect -4294 -3349 -4290 -3343
rect -4625 -3364 -4535 -3359
rect -4625 -3753 -4621 -3364
rect -4617 -3903 -4613 -3853
rect -4657 -3908 -4613 -3903
rect -4617 -4269 -4613 -3908
rect -4540 -3804 -4535 -3364
rect -4540 -4046 -4535 -3809
rect -4485 -3365 -4393 -3359
rect -4485 -3916 -4481 -3365
rect -4477 -4046 -4473 -4016
rect -4540 -4050 -4473 -4046
rect -6061 -4364 -6038 -4360
rect -6057 -4366 -6038 -4364
rect -6061 -4375 -6057 -4370
rect -6042 -4375 -6038 -4366
rect -6025 -4371 -6001 -4370
rect -6025 -4375 -6009 -4371
rect -6005 -4375 -6001 -4371
rect -6025 -4377 -6001 -4375
rect -6019 -4382 -6015 -4377
rect -6050 -4403 -6046 -4395
rect -6050 -4407 -6038 -4403
rect -6042 -4409 -6038 -4407
rect -6011 -4409 -6007 -4402
rect -5990 -4409 -5984 -4407
rect -6208 -4414 -6049 -4410
rect -6042 -4413 -6018 -4409
rect -6011 -4413 -5984 -4409
rect -6219 -4418 -6060 -4417
rect -6213 -4421 -6060 -4418
rect -6042 -4424 -6038 -4413
rect -6011 -4416 -6007 -4413
rect -6019 -4430 -6015 -4426
rect -6025 -4431 -6000 -4430
rect -6025 -4435 -6005 -4431
rect -6025 -4436 -6000 -4435
rect -6061 -4448 -6057 -4444
rect -6061 -4452 -6045 -4448
rect -6060 -4473 -6037 -4469
rect -6056 -4475 -6037 -4473
rect -6060 -4484 -6056 -4479
rect -6041 -4484 -6037 -4475
rect -6024 -4480 -6000 -4479
rect -6024 -4484 -6008 -4480
rect -6004 -4484 -6000 -4480
rect -6024 -4486 -6000 -4484
rect -6018 -4491 -6014 -4486
rect -6049 -4512 -6045 -4504
rect -6049 -4516 -6037 -4512
rect -6041 -4518 -6037 -4516
rect -6010 -4518 -6006 -4511
rect -5996 -4518 -5991 -4440
rect -6115 -4523 -6048 -4519
rect -6041 -4522 -6017 -4518
rect -6010 -4522 -5991 -4518
rect -6121 -4528 -6059 -4526
rect -6114 -4530 -6059 -4528
rect -6041 -4533 -6037 -4522
rect -6010 -4525 -6006 -4522
rect -6018 -4539 -6014 -4535
rect -6024 -4540 -5999 -4539
rect -6024 -4544 -6004 -4540
rect -6024 -4545 -5999 -4544
rect -6060 -4557 -6056 -4553
rect -6060 -4561 -6044 -4557
rect -6057 -4601 -6034 -4597
rect -6053 -4603 -6034 -4601
rect -6057 -4612 -6053 -4607
rect -6038 -4612 -6034 -4603
rect -6021 -4608 -5997 -4607
rect -6021 -4612 -6005 -4608
rect -6001 -4612 -5997 -4608
rect -6021 -4614 -5997 -4612
rect -6015 -4619 -6011 -4614
rect -6046 -4640 -6042 -4632
rect -6046 -4644 -6034 -4640
rect -6038 -4646 -6034 -4644
rect -6007 -4646 -6003 -4639
rect -5979 -4646 -5972 -4511
rect -6130 -4651 -6045 -4647
rect -6038 -4650 -6014 -4646
rect -6007 -4650 -5972 -4646
rect -6136 -4655 -6056 -4654
rect -6136 -4658 -6134 -4655
rect -6128 -4658 -6056 -4655
rect -6038 -4661 -6034 -4650
rect -6007 -4653 -6003 -4650
rect -6015 -4667 -6011 -4663
rect -6021 -4668 -5996 -4667
rect -6021 -4672 -6001 -4668
rect -6021 -4673 -5996 -4672
rect -6057 -4685 -6053 -4681
rect -6057 -4689 -6041 -4685
rect -6055 -4721 -6032 -4717
rect -6051 -4723 -6032 -4721
rect -6055 -4732 -6051 -4727
rect -6036 -4732 -6032 -4723
rect -6019 -4728 -5995 -4727
rect -6019 -4732 -6003 -4728
rect -5999 -4732 -5995 -4728
rect -6019 -4734 -5995 -4732
rect -6013 -4739 -6009 -4734
rect -6044 -4760 -6040 -4752
rect -6044 -4764 -6032 -4760
rect -6036 -4766 -6032 -4764
rect -6005 -4766 -6001 -4759
rect -5956 -4766 -5951 -4610
rect -6122 -4771 -6043 -4767
rect -6036 -4770 -6012 -4766
rect -6005 -4770 -5951 -4766
rect -6128 -4776 -6054 -4774
rect -6122 -4778 -6054 -4776
rect -6036 -4781 -6032 -4770
rect -6005 -4773 -6001 -4770
rect -6013 -4787 -6009 -4783
rect -6019 -4788 -5994 -4787
rect -6019 -4792 -5999 -4788
rect -6019 -4793 -5994 -4792
rect -6055 -4805 -6051 -4801
rect -6055 -4809 -6039 -4805
rect -6053 -4862 -6030 -4858
rect -6049 -4864 -6030 -4862
rect -6053 -4873 -6049 -4868
rect -6034 -4873 -6030 -4864
rect -6017 -4869 -5993 -4868
rect -6017 -4873 -6001 -4869
rect -5997 -4873 -5993 -4869
rect -6017 -4875 -5993 -4873
rect -6011 -4880 -6007 -4875
rect -6042 -4901 -6038 -4893
rect -6042 -4905 -6030 -4901
rect -6034 -4907 -6030 -4905
rect -6003 -4907 -5999 -4900
rect -5937 -4907 -5932 -4669
rect -5078 -4717 -5074 -4269
rect -4914 -4291 -4910 -4269
rect -4906 -4717 -4902 -4391
rect -4740 -4324 -4736 -4269
rect -4732 -4717 -4728 -4424
rect -4616 -4395 -4612 -4269
rect -4608 -4717 -4604 -4495
rect -4477 -4494 -4473 -4050
rect -4398 -3956 -4393 -3365
rect -4286 -3398 -4282 -3389
rect -4286 -3403 -4285 -3398
rect -4286 -3407 -4282 -3403
rect -4294 -3437 -4290 -3427
rect -4293 -3470 -4289 -3467
rect -4299 -3474 -4298 -3470
rect -4294 -3474 -4289 -3470
rect -4293 -3480 -4289 -3474
rect -4285 -3530 -4281 -3520
rect -4285 -3535 -4284 -3530
rect -4285 -3538 -4281 -3535
rect -4293 -3568 -4289 -3558
rect -4293 -3601 -4289 -3598
rect -4299 -3605 -4298 -3601
rect -4294 -3605 -4289 -3601
rect -4293 -3611 -4289 -3605
rect -4285 -3660 -4281 -3651
rect -4285 -3665 -4284 -3660
rect -4285 -3669 -4281 -3665
rect -4293 -3699 -4289 -3689
rect -4294 -3744 -4290 -3741
rect -4300 -3748 -4299 -3744
rect -4295 -3748 -4290 -3744
rect -4294 -3754 -4290 -3748
rect -4286 -3803 -4282 -3794
rect -4286 -3808 -4285 -3803
rect -4286 -3812 -4282 -3808
rect -4294 -3842 -4290 -3832
rect -4209 -3853 -4204 -2947
rect -4148 -3710 -4143 -2902
rect -4046 -3582 -4041 -2813
rect -3944 -3452 -3939 -2752
rect -3891 -3278 -3886 -2658
rect -3734 -3187 -3706 -3184
rect -3733 -3193 -3730 -3187
rect -3709 -3188 -3706 -3187
rect -3709 -3191 -3638 -3188
rect -3756 -3215 -3747 -3214
rect -3752 -3217 -3747 -3215
rect -3742 -3216 -3732 -3213
rect -3724 -3213 -3721 -3205
rect -3694 -3197 -3691 -3191
rect -3675 -3197 -3672 -3191
rect -3724 -3216 -3703 -3213
rect -3724 -3219 -3721 -3216
rect -3733 -3229 -3730 -3225
rect -3739 -3231 -3715 -3229
rect -3739 -3232 -3721 -3231
rect -3716 -3232 -3715 -3231
rect -3706 -3239 -3703 -3216
rect -3665 -3197 -3645 -3194
rect -3665 -3203 -3662 -3197
rect -3648 -3203 -3645 -3197
rect -3684 -3224 -3681 -3221
rect -3684 -3227 -3666 -3224
rect -3656 -3234 -3653 -3227
rect -3656 -3237 -3639 -3234
rect -3734 -3240 -3715 -3239
rect -3739 -3242 -3715 -3240
rect -3706 -3242 -3663 -3239
rect -3733 -3248 -3730 -3242
rect -3642 -3249 -3639 -3237
rect -3677 -3253 -3652 -3250
rect -3642 -3253 -3518 -3249
rect -3677 -3255 -3674 -3253
rect -3784 -3271 -3747 -3268
rect -3742 -3271 -3732 -3268
rect -3724 -3268 -3721 -3260
rect -3712 -3258 -3674 -3255
rect -3642 -3256 -3639 -3253
rect -3712 -3268 -3709 -3258
rect -3671 -3259 -3639 -3256
rect -3671 -3262 -3668 -3259
rect -3724 -3271 -3709 -3268
rect -3724 -3274 -3721 -3271
rect -3891 -3284 -3806 -3278
rect -3672 -3265 -3666 -3262
rect -3733 -3284 -3730 -3280
rect -3712 -3281 -3707 -3278
rect -3694 -3278 -3691 -3274
rect -3647 -3278 -3644 -3274
rect -3702 -3281 -3638 -3278
rect -3712 -3284 -3709 -3281
rect -3739 -3287 -3709 -3284
rect -3633 -3292 -3629 -3253
rect -3803 -3371 -3775 -3368
rect -3802 -3377 -3799 -3371
rect -3778 -3372 -3775 -3371
rect -3778 -3375 -3707 -3372
rect -3829 -3401 -3816 -3398
rect -3811 -3400 -3801 -3397
rect -3793 -3397 -3790 -3389
rect -3763 -3381 -3760 -3375
rect -3744 -3381 -3741 -3375
rect -3793 -3400 -3772 -3397
rect -3793 -3403 -3790 -3400
rect -3802 -3413 -3799 -3409
rect -3808 -3415 -3784 -3413
rect -3808 -3416 -3790 -3415
rect -3785 -3416 -3784 -3415
rect -3775 -3423 -3772 -3400
rect -3734 -3381 -3714 -3378
rect -3734 -3387 -3731 -3381
rect -3717 -3387 -3714 -3381
rect -3753 -3408 -3750 -3405
rect -3753 -3411 -3735 -3408
rect -3725 -3418 -3722 -3411
rect -3725 -3421 -3708 -3418
rect -3803 -3424 -3784 -3423
rect -3808 -3426 -3784 -3424
rect -3775 -3426 -3732 -3423
rect -3802 -3432 -3799 -3426
rect -3711 -3432 -3708 -3421
rect -3711 -3433 -3698 -3432
rect -3746 -3437 -3721 -3434
rect -3711 -3436 -3595 -3433
rect -3746 -3439 -3743 -3437
rect -3944 -3455 -3816 -3452
rect -3811 -3455 -3801 -3452
rect -3793 -3452 -3790 -3444
rect -3781 -3442 -3743 -3439
rect -3711 -3440 -3708 -3436
rect -3781 -3452 -3778 -3442
rect -3740 -3443 -3708 -3440
rect -3702 -3437 -3595 -3436
rect -3740 -3446 -3737 -3443
rect -3793 -3455 -3778 -3452
rect -3793 -3458 -3790 -3455
rect -3741 -3449 -3735 -3446
rect -3802 -3468 -3799 -3464
rect -3781 -3465 -3776 -3462
rect -3763 -3462 -3760 -3458
rect -3716 -3462 -3713 -3458
rect -3771 -3465 -3707 -3462
rect -3781 -3468 -3778 -3465
rect -3808 -3471 -3778 -3468
rect -3702 -3476 -3698 -3437
rect -3808 -3501 -3780 -3498
rect -3807 -3507 -3804 -3501
rect -3783 -3502 -3780 -3501
rect -3783 -3505 -3712 -3502
rect -3831 -3530 -3821 -3528
rect -3826 -3531 -3821 -3530
rect -3816 -3530 -3806 -3527
rect -3798 -3527 -3795 -3519
rect -3768 -3511 -3765 -3505
rect -3749 -3511 -3746 -3505
rect -3798 -3530 -3777 -3527
rect -3798 -3533 -3795 -3530
rect -3807 -3543 -3804 -3539
rect -3813 -3545 -3789 -3543
rect -3813 -3546 -3795 -3545
rect -3790 -3546 -3789 -3545
rect -3780 -3553 -3777 -3530
rect -3739 -3511 -3719 -3508
rect -3739 -3517 -3736 -3511
rect -3722 -3517 -3719 -3511
rect -3758 -3538 -3755 -3535
rect -3758 -3541 -3740 -3538
rect -3730 -3548 -3727 -3541
rect -3730 -3551 -3713 -3548
rect -3808 -3554 -3789 -3553
rect -3813 -3556 -3789 -3554
rect -3780 -3556 -3737 -3553
rect -3807 -3562 -3804 -3556
rect -3716 -3562 -3713 -3551
rect -3751 -3567 -3726 -3564
rect -3716 -3564 -3703 -3562
rect -3716 -3566 -3595 -3564
rect -3751 -3569 -3748 -3567
rect -4046 -3585 -3821 -3582
rect -3816 -3585 -3806 -3582
rect -3798 -3582 -3795 -3574
rect -3786 -3572 -3748 -3569
rect -3716 -3570 -3713 -3566
rect -3786 -3582 -3783 -3572
rect -3745 -3573 -3713 -3570
rect -3707 -3568 -3595 -3566
rect -3745 -3576 -3742 -3573
rect -3798 -3585 -3783 -3582
rect -3798 -3588 -3795 -3585
rect -3746 -3579 -3740 -3576
rect -3807 -3598 -3804 -3594
rect -3786 -3595 -3781 -3592
rect -3768 -3592 -3765 -3588
rect -3721 -3592 -3718 -3588
rect -3776 -3595 -3712 -3592
rect -3786 -3598 -3783 -3595
rect -3813 -3601 -3783 -3598
rect -3707 -3606 -3703 -3568
rect -3804 -3629 -3776 -3626
rect -3803 -3635 -3800 -3629
rect -3779 -3630 -3776 -3629
rect -3779 -3633 -3708 -3630
rect -3829 -3659 -3817 -3656
rect -3829 -3660 -3824 -3659
rect -3812 -3658 -3802 -3655
rect -3794 -3655 -3791 -3647
rect -3764 -3639 -3761 -3633
rect -3745 -3639 -3742 -3633
rect -3794 -3658 -3773 -3655
rect -3794 -3661 -3791 -3658
rect -3803 -3671 -3800 -3667
rect -3809 -3673 -3785 -3671
rect -3809 -3674 -3791 -3673
rect -3786 -3674 -3785 -3673
rect -3776 -3681 -3773 -3658
rect -3735 -3639 -3715 -3636
rect -3735 -3645 -3732 -3639
rect -3718 -3645 -3715 -3639
rect -3754 -3666 -3751 -3663
rect -3754 -3669 -3736 -3666
rect -3726 -3676 -3723 -3669
rect -3726 -3679 -3709 -3676
rect -3804 -3682 -3785 -3681
rect -3809 -3684 -3785 -3682
rect -3776 -3684 -3733 -3681
rect -3803 -3690 -3800 -3684
rect -3712 -3690 -3709 -3679
rect -3747 -3695 -3722 -3692
rect -3712 -3694 -3699 -3690
rect -3747 -3697 -3744 -3695
rect -4148 -3713 -3817 -3710
rect -3812 -3713 -3802 -3710
rect -3794 -3710 -3791 -3702
rect -3782 -3700 -3744 -3697
rect -3712 -3698 -3709 -3694
rect -3782 -3710 -3779 -3700
rect -3741 -3701 -3709 -3698
rect -3703 -3698 -3595 -3694
rect -3741 -3704 -3738 -3701
rect -3794 -3713 -3779 -3710
rect -3794 -3716 -3791 -3713
rect -3742 -3707 -3736 -3704
rect -3803 -3726 -3800 -3722
rect -3782 -3723 -3777 -3720
rect -3764 -3720 -3761 -3716
rect -3717 -3720 -3714 -3716
rect -3772 -3723 -3708 -3720
rect -3782 -3726 -3779 -3723
rect -3809 -3729 -3779 -3726
rect -3703 -3734 -3699 -3698
rect -3803 -3772 -3775 -3769
rect -3802 -3778 -3799 -3772
rect -3778 -3773 -3775 -3772
rect -3778 -3776 -3707 -3773
rect -3828 -3802 -3816 -3799
rect -3828 -3803 -3823 -3802
rect -3811 -3801 -3801 -3798
rect -3793 -3798 -3790 -3790
rect -3763 -3782 -3760 -3776
rect -3744 -3782 -3741 -3776
rect -3793 -3801 -3772 -3798
rect -3793 -3804 -3790 -3801
rect -3802 -3814 -3799 -3810
rect -3808 -3816 -3784 -3814
rect -3808 -3817 -3790 -3816
rect -3785 -3817 -3784 -3816
rect -3775 -3824 -3772 -3801
rect -3734 -3782 -3714 -3779
rect -3734 -3788 -3731 -3782
rect -3717 -3788 -3714 -3782
rect -3753 -3809 -3750 -3806
rect -3753 -3812 -3735 -3809
rect -3725 -3819 -3722 -3812
rect -3725 -3822 -3708 -3819
rect -3803 -3825 -3784 -3824
rect -3808 -3827 -3784 -3825
rect -3775 -3827 -3732 -3824
rect -3802 -3833 -3799 -3827
rect -3711 -3833 -3708 -3822
rect -3746 -3838 -3721 -3835
rect -3711 -3837 -3698 -3833
rect -3746 -3840 -3743 -3838
rect -4209 -3856 -3816 -3853
rect -3811 -3856 -3801 -3853
rect -3793 -3853 -3790 -3845
rect -3781 -3843 -3743 -3840
rect -3711 -3841 -3708 -3837
rect -3781 -3853 -3778 -3843
rect -3740 -3844 -3708 -3841
rect -3702 -3841 -3594 -3837
rect -3740 -3847 -3737 -3844
rect -3793 -3856 -3778 -3853
rect -3793 -3859 -3790 -3856
rect -3741 -3850 -3735 -3847
rect -3802 -3869 -3799 -3865
rect -3781 -3866 -3776 -3863
rect -3763 -3863 -3760 -3859
rect -3716 -3863 -3713 -3859
rect -3771 -3866 -3707 -3863
rect -3781 -3869 -3778 -3866
rect -3808 -3872 -3778 -3869
rect -3702 -3877 -3698 -3841
rect -4294 -3896 -4290 -3893
rect -4300 -3900 -4299 -3896
rect -4295 -3900 -4290 -3896
rect -4294 -3906 -4290 -3900
rect -4286 -3955 -4282 -3946
rect -4286 -3960 -4285 -3955
rect -4469 -4717 -4465 -4594
rect -4398 -4553 -4394 -3961
rect -4286 -3964 -4282 -3960
rect -4294 -3994 -4290 -3984
rect -5078 -4718 -4465 -4717
rect -4390 -4718 -4386 -4653
rect -5078 -4722 -4386 -4718
rect -5078 -4811 -5074 -4722
rect -5231 -4862 -5227 -4859
rect -5237 -4866 -5236 -4862
rect -5232 -4866 -5227 -4862
rect -6120 -4912 -6041 -4908
rect -6034 -4911 -6010 -4907
rect -6003 -4911 -5932 -4907
rect -5231 -4872 -5227 -4866
rect -6126 -4917 -6052 -4915
rect -6120 -4919 -6052 -4917
rect -6034 -4922 -6030 -4911
rect -6003 -4914 -5999 -4911
rect -5223 -4922 -5219 -4912
rect -5070 -4920 -5066 -4911
rect -6011 -4928 -6007 -4924
rect -5223 -4927 -5086 -4922
rect -6017 -4929 -5992 -4928
rect -6017 -4933 -5997 -4929
rect -5223 -4930 -5219 -4927
rect -6017 -4934 -5992 -4933
rect -6053 -4946 -6049 -4942
rect -6053 -4950 -6037 -4946
rect -5231 -4960 -5227 -4950
<< m2contact >>
rect -5882 -2602 -5877 -2595
rect -6293 -3476 -6288 -3471
rect -6091 -3477 -6086 -3472
rect -6276 -3532 -6271 -3527
rect -6091 -3531 -6086 -3526
rect -5977 -3515 -5972 -3510
rect -5984 -3604 -5979 -3599
rect -6186 -3650 -6181 -3645
rect -6098 -3649 -6093 -3644
rect -6185 -3704 -6180 -3699
rect -6098 -3703 -6093 -3698
rect -6176 -3794 -6171 -3789
rect -6095 -3793 -6090 -3788
rect -5765 -2666 -5760 -2659
rect -5765 -3515 -5760 -3510
rect -5708 -2752 -5703 -2745
rect -3944 -2752 -3939 -2746
rect -5708 -3604 -5703 -3599
rect -5616 -2813 -5611 -2806
rect -5882 -3783 -5877 -3778
rect -6183 -3848 -6178 -3843
rect -6095 -3847 -6090 -3842
rect -5981 -3838 -5976 -3833
rect -4046 -2813 -4041 -2807
rect -5616 -3838 -5611 -3833
rect -5487 -2902 -5482 -2895
rect -4148 -2902 -4143 -2895
rect -5985 -3869 -5980 -3864
rect -5487 -3869 -5482 -3864
rect -5327 -2947 -5322 -2942
rect -6179 -3942 -6174 -3937
rect -6099 -3941 -6094 -3936
rect -6179 -3996 -6174 -3991
rect -6099 -3995 -6094 -3990
rect -4209 -2947 -4204 -2942
rect -5115 -3290 -5108 -3284
rect -4942 -3291 -4937 -3285
rect -4997 -3404 -4992 -3399
rect -4768 -3291 -4762 -3285
rect -4644 -3292 -4639 -3286
rect -5960 -4032 -5955 -4027
rect -5327 -4032 -5322 -4027
rect -6154 -4158 -6149 -4153
rect -6074 -4157 -6069 -4152
rect -6154 -4212 -6149 -4207
rect -6074 -4211 -6069 -4206
rect -4814 -3535 -4809 -3530
rect -4657 -3666 -4652 -3661
rect -4504 -3295 -4499 -3289
rect -4540 -3809 -4535 -3804
rect -5990 -4407 -5984 -4402
rect -6213 -4414 -6208 -4409
rect -6219 -4423 -6213 -4418
rect -5996 -4440 -5991 -4435
rect -6121 -4523 -6115 -4518
rect -5979 -4511 -5972 -4506
rect -6121 -4534 -6114 -4528
rect -6136 -4651 -6130 -4646
rect -5956 -4610 -5951 -4605
rect -6134 -4660 -6128 -4655
rect -6128 -4771 -6122 -4765
rect -5937 -4669 -5932 -4664
rect -6128 -4781 -6122 -4776
rect -6126 -4912 -6120 -4906
rect -4285 -3403 -4280 -3398
rect -4284 -3535 -4279 -3530
rect -4284 -3665 -4279 -3660
rect -4285 -3808 -4280 -3803
rect -3758 -3220 -3752 -3215
rect -3747 -3218 -3742 -3213
rect -3789 -3273 -3784 -3268
rect -3747 -3272 -3742 -3267
rect -3806 -3284 -3799 -3278
rect -3834 -3403 -3829 -3398
rect -3816 -3402 -3811 -3397
rect -3816 -3456 -3811 -3451
rect -3831 -3535 -3826 -3530
rect -3821 -3532 -3816 -3527
rect -3821 -3586 -3816 -3581
rect -3817 -3660 -3812 -3655
rect -3829 -3665 -3824 -3660
rect -3817 -3714 -3812 -3709
rect -3816 -3803 -3811 -3798
rect -3828 -3808 -3823 -3803
rect -3816 -3857 -3811 -3852
rect -4398 -3961 -4393 -3956
rect -4285 -3960 -4280 -3955
rect -6126 -4922 -6120 -4917
rect -5086 -4927 -5081 -4922
<< pm12contact >>
rect -6035 -3494 -6030 -3489
rect -6026 -3495 -6021 -3490
rect -6042 -3666 -6037 -3661
rect -6033 -3667 -6028 -3662
rect -6039 -3810 -6034 -3805
rect -6030 -3811 -6025 -3806
rect -6043 -3958 -6038 -3953
rect -6034 -3959 -6029 -3954
rect -5237 -3045 -5232 -3040
rect -5104 -3290 -5098 -3284
rect -4932 -3291 -4926 -3285
rect -5095 -3515 -5090 -3510
rect -4758 -3291 -4752 -3285
rect -4634 -3292 -4628 -3286
rect -4923 -3604 -4918 -3599
rect -5087 -3783 -5082 -3778
rect -6018 -4174 -6013 -4169
rect -6009 -4175 -6004 -4170
rect -4749 -3838 -4744 -3833
rect -4494 -3295 -4488 -3289
rect -4625 -3869 -4620 -3864
rect -4485 -4032 -4480 -4027
rect -4914 -4407 -4909 -4402
rect -4740 -4440 -4735 -4435
rect -4616 -4511 -4611 -4506
rect -4294 -3404 -4289 -3399
rect -4293 -3535 -4288 -3530
rect -4293 -3666 -4288 -3661
rect -4294 -3809 -4289 -3804
rect -3691 -3235 -3686 -3230
rect -3682 -3236 -3677 -3231
rect -3760 -3419 -3755 -3414
rect -3751 -3420 -3746 -3415
rect -3765 -3549 -3760 -3544
rect -3756 -3550 -3751 -3545
rect -3761 -3677 -3756 -3672
rect -3752 -3678 -3747 -3673
rect -3760 -3820 -3755 -3815
rect -3751 -3821 -3746 -3816
rect -4294 -3961 -4289 -3956
rect -4477 -4610 -4472 -4605
rect -4398 -4669 -4393 -4664
rect -5231 -4927 -5226 -4922
rect -5078 -4927 -5073 -4922
<< metal2 >>
rect -5877 -2596 -4685 -2595
rect -5877 -2602 -3839 -2596
rect -5760 -2660 -4304 -2659
rect -5760 -2666 -3887 -2660
rect -5703 -2746 -4319 -2745
rect -5703 -2752 -3944 -2746
rect -5611 -2807 -4242 -2806
rect -5611 -2813 -4046 -2807
rect -5482 -2902 -4148 -2895
rect -5322 -2947 -4209 -2942
rect -5240 -3045 -5237 -3040
rect -3844 -3214 -3839 -2602
rect -3844 -3215 -3756 -3214
rect -3844 -3220 -3758 -3215
rect -3746 -3224 -3743 -3218
rect -3746 -3227 -3709 -3224
rect -3712 -3230 -3709 -3227
rect -3712 -3233 -3691 -3230
rect -3682 -3246 -3679 -3236
rect -3745 -3249 -3679 -3246
rect -3745 -3267 -3742 -3249
rect -3789 -3278 -3784 -3273
rect -3799 -3284 -3784 -3278
rect -5108 -3290 -5104 -3284
rect -4937 -3291 -4932 -3285
rect -4762 -3291 -4758 -3285
rect -4639 -3292 -4634 -3286
rect -4499 -3295 -4494 -3289
rect -4992 -3404 -4294 -3399
rect -4280 -3403 -3834 -3398
rect -3815 -3408 -3812 -3402
rect -3815 -3411 -3778 -3408
rect -3781 -3414 -3778 -3411
rect -3781 -3417 -3760 -3414
rect -3751 -3430 -3748 -3420
rect -3814 -3433 -3748 -3430
rect -3814 -3451 -3811 -3433
rect -6385 -3476 -6293 -3471
rect -6090 -3483 -6087 -3477
rect -6090 -3486 -6053 -3483
rect -6056 -3489 -6053 -3486
rect -6056 -3492 -6035 -3489
rect -6026 -3505 -6023 -3495
rect -6089 -3508 -6023 -3505
rect -6089 -3526 -6086 -3508
rect -5972 -3515 -5765 -3510
rect -5760 -3515 -5095 -3510
rect -6385 -3532 -6276 -3527
rect -4809 -3535 -4293 -3530
rect -4279 -3535 -3831 -3530
rect -3820 -3538 -3817 -3532
rect -3820 -3541 -3783 -3538
rect -3786 -3544 -3783 -3541
rect -3786 -3547 -3765 -3544
rect -3756 -3560 -3753 -3550
rect -3819 -3563 -3753 -3560
rect -3819 -3581 -3816 -3563
rect -5979 -3604 -5708 -3599
rect -5703 -3604 -4923 -3599
rect -6385 -3650 -6186 -3645
rect -6097 -3655 -6094 -3649
rect -6097 -3658 -6060 -3655
rect -6063 -3661 -6060 -3658
rect -6063 -3664 -6042 -3661
rect -4652 -3666 -4293 -3661
rect -4279 -3665 -3829 -3660
rect -3816 -3666 -3813 -3660
rect -6033 -3677 -6030 -3667
rect -3816 -3669 -3779 -3666
rect -3782 -3672 -3779 -3669
rect -6096 -3680 -6030 -3677
rect -6096 -3698 -6093 -3680
rect -3782 -3675 -3761 -3672
rect -3752 -3688 -3749 -3678
rect -6385 -3704 -6185 -3699
rect -3815 -3691 -3749 -3688
rect -3815 -3709 -3812 -3691
rect -5877 -3783 -5087 -3778
rect -6385 -3794 -6176 -3789
rect -6094 -3799 -6091 -3793
rect -6094 -3802 -6057 -3799
rect -6060 -3805 -6057 -3802
rect -6060 -3808 -6039 -3805
rect -4535 -3809 -4294 -3804
rect -4280 -3808 -3828 -3803
rect -3815 -3809 -3812 -3803
rect -6030 -3821 -6027 -3811
rect -3815 -3812 -3778 -3809
rect -3781 -3815 -3778 -3812
rect -6093 -3824 -6027 -3821
rect -6093 -3842 -6090 -3824
rect -3781 -3818 -3760 -3815
rect -3751 -3831 -3748 -3821
rect -5976 -3838 -5616 -3833
rect -5611 -3838 -4749 -3833
rect -3814 -3834 -3748 -3831
rect -6385 -3848 -6183 -3843
rect -3814 -3852 -3811 -3834
rect -5980 -3869 -5487 -3864
rect -5482 -3869 -4625 -3864
rect -6385 -3942 -6179 -3937
rect -6098 -3947 -6095 -3941
rect -6098 -3950 -6061 -3947
rect -6064 -3953 -6061 -3950
rect -6064 -3956 -6043 -3953
rect -6034 -3969 -6031 -3959
rect -4393 -3961 -4294 -3956
rect -4280 -3960 -3605 -3955
rect -6097 -3972 -6031 -3969
rect -6097 -3990 -6094 -3972
rect -6385 -3996 -6179 -3991
rect -5955 -4032 -5327 -4027
rect -5322 -4032 -4485 -4027
rect -6360 -4158 -6154 -4153
rect -6073 -4163 -6070 -4157
rect -6073 -4166 -6036 -4163
rect -6039 -4169 -6036 -4166
rect -6039 -4172 -6018 -4169
rect -6009 -4185 -6006 -4175
rect -6072 -4188 -6006 -4185
rect -6072 -4206 -6069 -4188
rect -6360 -4212 -6154 -4207
rect -5984 -4407 -4914 -4402
rect -6384 -4413 -6213 -4409
rect -6384 -4418 -6221 -4417
rect -6384 -4422 -6219 -4418
rect -6219 -4425 -6213 -4423
rect -5991 -4440 -4740 -4435
rect -5972 -4511 -4616 -4506
rect -6146 -4522 -6121 -4518
rect -6384 -4523 -6121 -4522
rect -6384 -4526 -6140 -4523
rect -6384 -4534 -6121 -4530
rect -6384 -4535 -6114 -4534
rect -5951 -4610 -4477 -4605
rect -6158 -4647 -6136 -4646
rect -6384 -4651 -6136 -4647
rect -6384 -4660 -6134 -4655
rect -6128 -4660 -6127 -4655
rect -5932 -4669 -4398 -4664
rect -6156 -4769 -6128 -4765
rect -6384 -4771 -6128 -4769
rect -6122 -4771 -6121 -4767
rect -6384 -4772 -6121 -4771
rect -6384 -4773 -6154 -4772
rect -6384 -4781 -6128 -4777
rect -6122 -4781 -6121 -4777
rect -6384 -4782 -6121 -4781
rect -6154 -4910 -6126 -4906
rect -6382 -4912 -6126 -4910
rect -6120 -4912 -6119 -4908
rect -6382 -4913 -6119 -4912
rect -6382 -4914 -6152 -4913
rect -6382 -4922 -6126 -4918
rect -6120 -4922 -6119 -4918
rect -6382 -4923 -6119 -4922
rect -5241 -4927 -5231 -4922
rect -5081 -4927 -5078 -4922
<< m123contact >>
rect -3739 -3187 -3734 -3182
rect -3739 -3240 -3734 -3235
rect -3721 -3236 -3716 -3231
rect -3707 -3281 -3702 -3276
rect -3808 -3371 -3803 -3366
rect -3808 -3424 -3803 -3419
rect -3790 -3420 -3785 -3415
rect -6083 -3446 -6078 -3441
rect -3776 -3465 -3771 -3460
rect -6083 -3499 -6078 -3494
rect -6065 -3495 -6060 -3490
rect -3813 -3501 -3808 -3496
rect -6051 -3540 -6046 -3535
rect -3813 -3554 -3808 -3549
rect -3795 -3550 -3790 -3545
rect -3781 -3595 -3776 -3590
rect -6090 -3618 -6085 -3613
rect -3809 -3629 -3804 -3624
rect -6090 -3671 -6085 -3666
rect -6072 -3667 -6067 -3662
rect -3809 -3682 -3804 -3677
rect -3791 -3678 -3786 -3673
rect -6058 -3712 -6053 -3707
rect -3777 -3723 -3772 -3718
rect -6087 -3762 -6082 -3757
rect -3808 -3772 -3803 -3767
rect -6087 -3815 -6082 -3810
rect -6069 -3811 -6064 -3806
rect -3808 -3825 -3803 -3820
rect -3790 -3821 -3785 -3816
rect -6055 -3856 -6050 -3851
rect -3776 -3866 -3771 -3861
rect -6091 -3910 -6086 -3905
rect -6091 -3963 -6086 -3958
rect -6073 -3959 -6068 -3954
rect -6059 -4004 -6054 -3999
rect -6066 -4126 -6061 -4121
rect -6066 -4179 -6061 -4174
rect -6048 -4175 -6043 -4170
rect -6034 -4220 -6029 -4215
<< metal3 >>
rect -3739 -3235 -3736 -3187
rect -3716 -3236 -3704 -3233
rect -3707 -3276 -3704 -3236
rect -3808 -3419 -3805 -3371
rect -3785 -3420 -3773 -3417
rect -6083 -3494 -6080 -3446
rect -3776 -3460 -3773 -3420
rect -6060 -3495 -6048 -3492
rect -6051 -3535 -6048 -3495
rect -3813 -3549 -3810 -3501
rect -3790 -3550 -3778 -3547
rect -3781 -3590 -3778 -3550
rect -6090 -3666 -6087 -3618
rect -6067 -3667 -6055 -3664
rect -6058 -3707 -6055 -3667
rect -3809 -3677 -3806 -3629
rect -3786 -3678 -3774 -3675
rect -3777 -3718 -3774 -3678
rect -6087 -3810 -6084 -3762
rect -6064 -3811 -6052 -3808
rect -6055 -3851 -6052 -3811
rect -3808 -3820 -3805 -3772
rect -3785 -3821 -3773 -3818
rect -3776 -3861 -3773 -3821
rect -6091 -3958 -6088 -3910
rect -6068 -3959 -6056 -3956
rect -6059 -3999 -6056 -3959
rect -6066 -4174 -6063 -4126
rect -6043 -4175 -6031 -4172
rect -6034 -4215 -6031 -4175
<< labels >>
rlabel metal2 -3610 -3958 -3609 -3957 1 cout
rlabel metal1 -4294 -3994 -4290 -3990 1 gnd!
rlabel metal1 -4294 -3896 -4290 -3893 1 vdd!
rlabel metal1 -5958 -4033 -5958 -4031 1 prop_5
rlabel metal1 -3721 -3287 -3717 -3284 1 gnd
rlabel metal1 -3671 -3281 -3668 -3279 1 gnd
rlabel metal1 -3723 -3231 -3722 -3229 1 gnd
rlabel metal1 -3727 -3187 -3724 -3185 5 vdd
rlabel metal1 -3726 -3241 -3723 -3239 1 vdd
rlabel metal1 -3630 -3250 -3630 -3250 1 s1
rlabel m2contact -3788 -3269 -3788 -3269 1 prop_1
rlabel metal1 -3701 -3836 -3699 -3834 1 s5
rlabel metal1 -3817 -3854 -3815 -3854 1 prop_5
rlabel metal1 -3795 -3826 -3792 -3824 1 vdd
rlabel metal1 -3796 -3772 -3793 -3770 5 vdd
rlabel metal1 -3792 -3816 -3791 -3814 1 gnd
rlabel metal1 -3740 -3866 -3737 -3864 1 gnd
rlabel metal1 -3790 -3872 -3786 -3869 1 gnd
rlabel metal1 -4390 -4662 -4386 -4657 7 clock_car0
rlabel m2contact -6126 -4922 -6120 -4917 1 q_b5
rlabel m2contact -6126 -4912 -6120 -4906 1 q_a5
rlabel metal1 -6013 -4873 -6013 -4873 5 vdd
rlabel metal1 -6010 -4930 -6010 -4930 1 gnd
rlabel metal1 -6042 -4948 -6042 -4948 1 gnd
rlabel metal1 -6043 -4861 -6043 -4861 5 vdd
rlabel metal1 -4493 -3207 -4489 -3202 5 vdd!
rlabel metal2 -4504 -3295 -4499 -3289 1 clock_in
rlabel metal1 -4469 -4603 -4465 -4598 7 clock_car0
rlabel metal2 -4485 -4610 -4481 -4605 1 gen_4
rlabel metal1 -4477 -4491 -4473 -4486 1 pdr4
rlabel metal1 -4477 -4046 -4473 -4016 1 pdr4
rlabel metal2 -4500 -4032 -4485 -4027 1 prop_5
rlabel metal1 -4485 -3916 -4481 -3899 1 pdr5
rlabel m2contact -6154 -4212 -6149 -4207 1 q_b5
rlabel m2contact -6154 -4158 -6149 -4153 1 q_a5
rlabel metal1 -6053 -4180 -6050 -4178 1 vdd
rlabel metal1 -6054 -4126 -6051 -4124 5 vdd
rlabel metal1 -6050 -4170 -6049 -4168 1 gnd
rlabel metal1 -5998 -4220 -5995 -4218 1 gnd
rlabel metal1 -6048 -4226 -6044 -4223 1 gnd
rlabel m2contact -6127 -4769 -6127 -4769 3 q_a4
rlabel m2contact -6212 -4412 -6212 -4412 3 q_a1
rlabel metal1 -6127 -4775 -6127 -4775 3 q_b4
rlabel m2contact -6119 -4529 -6119 -4529 1 q_b2
rlabel m2contact -6119 -4522 -6119 -4522 1 q_a2
rlabel metal1 -5997 -4768 -5997 -4768 1 gen_4
rlabel metal1 -6015 -4732 -6015 -4732 5 vdd
rlabel metal1 -6012 -4789 -6012 -4789 1 gnd
rlabel metal1 -6044 -4807 -6044 -4807 1 gnd
rlabel metal1 -6045 -4720 -6045 -4720 5 vdd
rlabel metal1 -5974 -4648 -5974 -4648 1 gen_3
rlabel metal1 -6017 -4612 -6017 -4612 5 vdd
rlabel metal1 -6014 -4669 -6014 -4669 1 gnd
rlabel metal1 -6046 -4687 -6046 -4687 1 gnd
rlabel metal1 -6047 -4600 -6047 -4600 5 vdd
rlabel metal1 -5992 -4520 -5992 -4520 1 gen_2
rlabel metal1 -6020 -4484 -6020 -4484 5 vdd
rlabel metal1 -6017 -4541 -6017 -4541 1 gnd
rlabel metal1 -6049 -4559 -6049 -4559 1 gnd
rlabel metal1 -6050 -4472 -6050 -4472 5 vdd
rlabel metal1 -5985 -4412 -5985 -4412 1 gen_1
rlabel metal1 -6064 -4419 -6064 -4419 3 q_b1
rlabel metal1 -6021 -4375 -6021 -4375 5 vdd
rlabel metal1 -6018 -4432 -6018 -4432 1 gnd
rlabel metal1 -6050 -4450 -6050 -4450 1 gnd
rlabel metal1 -6051 -4363 -6051 -4363 5 vdd
rlabel metal1 -5070 -4920 -5066 -4916 1 gnd!
rlabel metal1 -5078 -4807 -5074 -4803 1 clock_car0
rlabel metal1 -4608 -4504 -4604 -4500 1 clock_car0
rlabel metal2 -4624 -4511 -4620 -4506 1 gen_3
rlabel metal1 -4616 -4392 -4612 -4387 1 pdr3
rlabel metal1 -4906 -4400 -4902 -4396 1 clock_car0
rlabel metal2 -4922 -4407 -4918 -4402 1 gen_1
rlabel metal1 -4914 -4288 -4910 -4283 1 pdr1
rlabel metal1 -4732 -4433 -4728 -4428 1 clock_car0
rlabel metal2 -4748 -4440 -4744 -4435 1 gen_2
rlabel metal1 -4740 -4321 -4736 -4316 1 pdr2
rlabel m2contact -6184 -3701 -6184 -3701 3 q_b2
rlabel m2contact -6178 -3939 -6178 -3939 1 q_a4
rlabel m2contact -6292 -3474 -6292 -3474 1 q_a1
rlabel m2contact -6275 -3528 -6275 -3528 1 q_b1
rlabel m2contact -6178 -3992 -6178 -3992 1 q_b4
rlabel m2contact -6185 -3646 -6185 -3646 3 q_a2
rlabel metal1 -5879 -3172 -5879 -3172 1 carry_0
rlabel metal1 -3943 -3454 -3943 -3454 1 prop_2
rlabel metal1 -3819 -3711 -3819 -3711 1 prop_4
rlabel metal1 -3701 -3692 -3701 -3692 1 s4
rlabel metal1 -3796 -3683 -3793 -3681 1 vdd
rlabel metal1 -3797 -3629 -3794 -3627 5 vdd
rlabel metal1 -3793 -3673 -3792 -3671 1 gnd
rlabel metal1 -3741 -3723 -3738 -3721 1 gnd
rlabel metal1 -3791 -3729 -3787 -3726 1 gnd
rlabel metal1 -3830 -3529 -3830 -3529 1 c2
rlabel metal1 -3795 -3601 -3791 -3598 1 gnd
rlabel metal1 -3745 -3595 -3742 -3593 1 gnd
rlabel metal1 -3797 -3545 -3796 -3543 1 gnd
rlabel metal1 -3801 -3501 -3798 -3499 5 vdd
rlabel metal1 -3800 -3555 -3797 -3553 1 vdd
rlabel metal1 -3823 -3584 -3823 -3584 1 prop_3
rlabel metal1 -3704 -3564 -3704 -3564 1 s3
rlabel metal1 -3699 -3435 -3699 -3435 7 s2
rlabel metal1 -3817 -3400 -3817 -3400 1 c1
rlabel metal1 -3795 -3425 -3792 -3423 1 vdd
rlabel metal1 -3796 -3371 -3793 -3369 5 vdd
rlabel metal1 -3792 -3415 -3791 -3413 1 gnd
rlabel metal1 -3740 -3465 -3737 -3463 1 gnd
rlabel metal1 -3790 -3471 -3786 -3468 1 gnd
rlabel metal1 -5982 -3878 -5982 -3878 1 prop_4
rlabel metal1 -6078 -3964 -6075 -3962 1 vdd
rlabel metal1 -6079 -3910 -6076 -3908 5 vdd
rlabel metal1 -6075 -3954 -6074 -3952 1 gnd
rlabel metal1 -6023 -4004 -6020 -4002 1 gnd
rlabel metal1 -6073 -4010 -6069 -4007 1 gnd
rlabel metal1 -5979 -3825 -5979 -3825 1 prop_3
rlabel metal1 -6096 -3844 -6096 -3844 1 q_b3
rlabel metal1 -6096 -3790 -6096 -3790 1 q_a3
rlabel metal1 -6074 -3816 -6071 -3814 1 vdd
rlabel metal1 -6075 -3762 -6072 -3760 5 vdd
rlabel metal1 -6071 -3806 -6070 -3804 1 gnd
rlabel metal1 -6019 -3856 -6016 -3854 1 gnd
rlabel metal1 -6069 -3862 -6065 -3859 1 gnd
rlabel metal1 -5982 -3680 -5982 -3680 1 prop_2
rlabel metal1 -6077 -3672 -6074 -3670 1 vdd
rlabel metal1 -6078 -3618 -6075 -3616 5 vdd
rlabel metal1 -6074 -3662 -6073 -3660 1 gnd
rlabel metal1 -6022 -3712 -6019 -3710 1 gnd
rlabel metal1 -6072 -3718 -6068 -3715 1 gnd
rlabel metal1 -5977 -3509 -5977 -3509 1 prop_1
rlabel metal1 -6070 -3500 -6067 -3498 1 vdd
rlabel metal1 -6071 -3446 -6068 -3444 5 vdd
rlabel metal1 -6067 -3490 -6066 -3488 1 gnd
rlabel metal1 -6015 -3540 -6012 -3538 1 gnd
rlabel metal1 -6065 -3546 -6061 -3543 1 gnd
rlabel metal1 -4285 -3809 -4282 -3804 1 c4
rlabel metal2 -4297 -3809 -4295 -3804 1 pdr4
rlabel metal1 -4294 -3842 -4290 -3838 1 gnd!
rlabel metal1 -4294 -3744 -4290 -3741 1 vdd!
rlabel metal2 -4657 -3666 -4655 -3661 1 pdr3
rlabel metal1 -4284 -3666 -4281 -3661 1 c3
rlabel metal1 -4293 -3699 -4289 -3695 1 gnd!
rlabel metal1 -4293 -3601 -4289 -3598 1 vdd!
rlabel metal1 -4293 -3471 -4289 -3467 1 vdd!
rlabel metal1 -4293 -3568 -4289 -3564 1 gnd!
rlabel metal2 -4296 -3535 -4294 -3530 1 pdr2
rlabel m2contact -4284 -3535 -4281 -3530 1 c2
rlabel metal2 -4997 -3404 -4995 -3399 1 pdr1
rlabel metal1 -4285 -3404 -4282 -3400 1 c1
rlabel metal1 -4294 -3437 -4290 -3433 1 gnd!
rlabel metal1 -4294 -3340 -4290 -3336 1 vdd!
rlabel metal1 -4617 -3862 -4613 -3858 1 pdr3
rlabel metal2 -4633 -3869 -4629 -3864 1 prop_4
rlabel metal1 -4625 -3749 -4621 -3745 1 pdr4
rlabel metal1 -4741 -3831 -4737 -3827 1 pdr2
rlabel metal2 -4757 -3838 -4753 -3833 1 prop_3
rlabel metal1 -4749 -3719 -4745 -3714 1 pdr3
rlabel metal1 -5087 -3664 -5083 -3659 1 prop1_car0
rlabel metal2 -5095 -3783 -5091 -3778 1 carry_0
rlabel metal1 -5079 -3776 -5075 -3771 1 clock_car0
rlabel metal1 -5087 -3508 -5083 -3503 1 prop1_car0
rlabel metal2 -5103 -3515 -5098 -3510 2 prop_1
rlabel metal1 -5095 -3396 -5091 -3391 1 pdr1
rlabel metal1 -4915 -3597 -4911 -3592 1 pdr1
rlabel metal2 -4931 -3604 -4926 -3599 1 prop_2
rlabel metal1 -4923 -3485 -4919 -3480 1 pdr2
rlabel metal1 -4633 -3204 -4629 -3199 5 vdd!
rlabel metal2 -4644 -3292 -4639 -3286 1 clock_in
rlabel metal1 -4625 -3283 -4621 -3279 1 pdr4
rlabel metal1 -4749 -3282 -4745 -3278 1 pdr3
rlabel metal2 -4768 -3291 -4762 -3285 1 clock_in
rlabel metal1 -4757 -3203 -4753 -3198 5 vdd!
rlabel metal1 -4931 -3203 -4927 -3198 5 vdd!
rlabel metal2 -4942 -3291 -4936 -3285 1 clock_in
rlabel metal1 -4923 -3282 -4919 -3278 1 pdr2
rlabel metal1 -5095 -3281 -5091 -3276 1 pdr1
rlabel metal2 -5114 -3290 -5108 -3284 2 clock_in
rlabel metal1 -5103 -3202 -5099 -3197 5 vdd!
rlabel metal1 -5228 -3045 -5225 -3041 1 clock_in
rlabel metal2 -5240 -3045 -5237 -3040 1 clk_org
rlabel metal1 -5237 -3078 -5233 -3074 1 gnd!
rlabel metal1 -5237 -2981 -5233 -2977 1 vdd!
rlabel metal1 -5996 -4910 -5994 -4908 1 gen_5
rlabel metal2 -4406 -4669 -4402 -4664 1 gen_5
rlabel metal2 -4297 -3961 -4295 -3956 1 pdr5
rlabel metal1 -4398 -4550 -4394 -4545 1 pdr5
rlabel metal1 -4485 -3286 -4481 -3282 1 pdr5
rlabel m2contact -6136 -4651 -6134 -4649 1 q_a3
rlabel metal1 -6061 -4658 -6059 -4656 1 q_b3
rlabel metal2 -5086 -4927 -5081 -4922 1 clock_in
rlabel metal1 -5222 -4927 -5219 -4923 1 clock_in
rlabel metal2 -5234 -4927 -5231 -4922 1 clk_org
rlabel metal1 -5231 -4960 -5227 -4956 1 gnd!
rlabel metal1 -5231 -4863 -5227 -4859 1 vdd!
<< end >>
