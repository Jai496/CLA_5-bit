magic
tech scmos
timestamp 1764616623
<< nwell >>
rect -143 66 -118 89
rect -100 66 -75 87
rect -58 66 -33 89
rect -2 69 55 94
rect 73 66 98 89
rect 116 66 141 87
rect 158 66 183 89
rect 214 69 271 94
<< ntransistor >>
rect -132 54 -130 58
rect -89 53 -87 57
rect -47 54 -45 58
rect 14 51 16 55
rect 35 51 37 55
rect 84 54 86 58
rect 127 53 129 57
rect 169 54 171 58
rect 230 51 232 55
rect 251 51 253 55
<< ptransistor >>
rect -132 73 -130 81
rect -89 73 -87 81
rect -47 73 -45 81
rect 14 76 16 84
rect 35 76 37 84
rect 84 73 86 81
rect 127 73 129 81
rect 169 73 171 81
rect 230 76 232 84
rect 251 76 253 84
<< ndiffusion >>
rect -133 54 -132 58
rect -130 54 -129 58
rect -90 53 -89 57
rect -87 53 -86 57
rect -48 54 -47 58
rect -45 54 -44 58
rect 13 51 14 55
rect 16 51 17 55
rect 34 51 35 55
rect 37 51 38 55
rect 83 54 84 58
rect 86 54 87 58
rect 126 53 127 57
rect 129 53 130 57
rect 168 54 169 58
rect 171 54 172 58
rect 229 51 230 55
rect 232 51 233 55
rect 250 51 251 55
rect 253 51 254 55
<< pdiffusion >>
rect -133 73 -132 81
rect -130 73 -129 81
rect -90 73 -89 81
rect -87 73 -86 81
rect -48 73 -47 81
rect -45 73 -44 81
rect 13 76 14 84
rect 16 76 17 84
rect 34 76 35 84
rect 37 76 38 84
rect 83 73 84 81
rect 86 73 87 81
rect 126 73 127 81
rect 129 73 130 81
rect 168 73 169 81
rect 171 73 172 81
rect 229 76 230 84
rect 232 76 233 84
rect 250 76 251 84
rect 253 76 254 84
<< ndcontact >>
rect -137 54 -133 58
rect -129 54 -125 58
rect -94 53 -90 57
rect -86 53 -82 57
rect -52 54 -48 58
rect -44 54 -40 58
rect 9 51 13 55
rect 17 51 21 55
rect 30 51 34 55
rect 38 51 42 55
rect 79 54 83 58
rect 87 54 91 58
rect 122 53 126 57
rect 130 53 134 57
rect 164 54 168 58
rect 172 54 176 58
rect 225 51 229 55
rect 233 51 237 55
rect 246 51 250 55
rect 254 51 258 55
<< pdcontact >>
rect -137 73 -133 81
rect -129 73 -125 81
rect -94 73 -90 81
rect -86 73 -82 81
rect -52 73 -48 81
rect -44 73 -40 81
rect 9 76 13 84
rect 17 76 21 84
rect 30 76 34 84
rect 38 76 42 84
rect 79 73 83 81
rect 87 73 91 81
rect 122 73 126 81
rect 130 73 134 81
rect 164 73 168 81
rect 172 73 176 81
rect 225 76 229 84
rect 233 76 237 84
rect 246 76 250 84
rect 254 76 258 84
<< polysilicon >>
rect -89 83 -87 100
rect 14 85 16 87
rect 35 84 37 103
rect 127 83 129 100
rect 230 85 232 87
rect 251 84 253 103
rect -132 58 -130 73
rect -89 66 -87 73
rect -89 57 -87 62
rect -47 58 -45 73
rect -132 51 -130 54
rect 14 55 16 76
rect 35 72 37 76
rect 84 58 86 73
rect 127 66 129 73
rect 35 55 37 58
rect -89 39 -87 53
rect -47 51 -45 54
rect 127 57 129 62
rect 169 58 171 73
rect 84 51 86 54
rect 230 55 232 76
rect 251 72 253 76
rect 251 55 253 58
rect 14 48 16 51
rect 35 35 37 51
rect 127 39 129 53
rect 169 51 171 54
rect 230 48 232 51
rect 251 35 253 51
<< polycontact >>
rect -93 96 -89 100
rect 31 99 35 103
rect 123 96 127 100
rect 247 99 251 103
rect -136 61 -132 65
rect -51 61 -47 65
rect 10 61 14 65
rect 80 61 84 65
rect -93 39 -89 43
rect 165 61 169 65
rect 226 61 230 65
rect 31 35 35 39
rect 123 39 127 43
rect 247 35 251 39
<< polypplus >>
rect -132 81 -130 84
rect 14 84 16 85
rect -89 81 -87 83
rect -47 81 -45 84
rect 84 81 86 84
rect 230 84 232 85
rect 127 81 129 83
rect 169 81 171 84
<< metal1 >>
rect -105 96 -93 100
rect 21 99 31 103
rect 111 96 123 100
rect 237 99 247 103
rect -143 85 -118 89
rect -58 85 -33 89
rect 9 88 34 92
rect -137 81 -133 85
rect -52 81 -48 85
rect 9 84 13 88
rect 30 84 34 88
rect -129 65 -125 73
rect -94 65 -90 73
rect -159 61 -136 65
rect -129 61 -90 65
rect -129 58 -125 61
rect -94 57 -90 61
rect -137 50 -133 54
rect 38 88 51 92
rect 38 84 42 88
rect 73 85 98 89
rect 158 85 183 89
rect 225 88 250 92
rect 79 81 83 85
rect 164 81 168 85
rect 225 84 229 88
rect 246 84 250 88
rect -86 65 -82 73
rect -44 65 -40 73
rect 17 65 21 76
rect 87 65 91 73
rect 122 65 126 73
rect -86 61 -51 65
rect -44 61 10 65
rect 17 61 80 65
rect 87 61 126 65
rect -86 57 -82 61
rect -44 58 -40 61
rect 17 55 21 61
rect 87 58 91 61
rect -52 50 -48 54
rect -143 47 -118 50
rect -58 47 -33 50
rect 9 46 13 51
rect 30 46 34 51
rect -107 39 -93 43
rect 9 42 34 46
rect 38 46 42 51
rect 122 57 126 61
rect 79 50 83 54
rect 254 88 267 92
rect 254 84 258 88
rect 130 65 134 73
rect 172 65 176 73
rect 233 65 237 76
rect 130 61 165 65
rect 172 61 226 65
rect 233 61 273 65
rect 130 57 134 61
rect 172 58 176 61
rect 233 55 237 61
rect 164 50 168 54
rect 73 47 98 50
rect 158 47 183 50
rect 225 46 229 51
rect 246 46 250 51
rect 38 42 51 46
rect 109 39 123 43
rect 225 42 250 46
rect 254 46 258 51
rect 254 42 267 46
rect -107 36 -103 39
rect 22 35 31 39
rect 238 35 247 39
<< labels >>
rlabel metal1 21 100 22 102 5 CLK
rlabel metal1 22 35 23 39 1 CLK_bar
rlabel metal1 49 89 50 91 1 vdd!
rlabel metal1 49 43 50 45 1 gnd!
rlabel metal1 -143 85 -118 89 1 vdd!
rlabel metal1 -143 47 -118 50 1 gnd!
rlabel metal1 -43 48 -42 49 1 gnd!
rlabel metal1 -48 87 -47 88 1 vdd!
rlabel metal1 265 89 266 91 1 vdd!
rlabel metal1 265 43 266 45 1 gnd!
rlabel metal1 73 85 98 89 1 vdd!
rlabel metal1 73 47 98 50 1 gnd!
rlabel metal1 159 62 160 63 1 storage
rlabel metal1 184 62 186 63 1 storage_bar
rlabel metal1 99 63 101 64 1 node1
rlabel metal1 233 43 235 45 1 storage_bar_gnd
rlabel metal1 232 89 234 91 1 storage_bar_vdd
rlabel metal1 173 48 174 49 1 gnd!
rlabel metal1 168 87 169 88 1 vdd!
rlabel metal1 238 35 239 39 1 CLK
rlabel metal1 237 100 238 102 5 CLK_bar
rlabel metal1 -117 63 -115 64 1 neg_node1
rlabel metal1 -57 62 -56 63 1 neg_storage
rlabel metal1 -32 62 -30 63 1 neg_storage_bar
rlabel metal1 17 43 19 45 1 neg_storage_bar_gnd
rlabel metal1 16 89 18 91 1 neg_storage_bar_vdd
rlabel metal1 -158 62 -157 63 3 FF_in
rlabel metal1 268 62 270 64 7 FF_out
rlabel metal1 111 96 114 100 5 clock_org
rlabel metal1 109 39 112 43 1 clock_in
rlabel metal1 -105 96 -102 100 5 clock_org
rlabel metal1 -107 39 -103 43 1 clock_in
<< end >>
